magic
tech sky130A
timestamp 1654986623
<< metal1 >>
rect 1300 7000 1400 7100
rect 1400 7100 1400 7100
rect 1500 7100 1500 7100
rect 1600 7100 1600 7100
rect 1700 7100 1700 7100
rect 1300 7100 1300 7200
rect 1700 7100 1800 7200
rect 1400 7200 1400 7200
rect 1800 7200 1800 7200
rect 1500 7200 1500 7200
rect 1900 7200 1900 7200
rect 1600 7200 1600 7200
rect 2000 7200 2000 7200
rect 1600 7200 1700 7200
rect 1700 7200 1700 7300
rect 1800 7300 1800 7300
rect 1800 7300 1800 7300
rect 1700 7300 1700 7300
rect 1700 7300 1700 7300
rect 1600 7300 1600 7400
rect 1900 7300 1900 7400
rect 1500 7400 1500 7400
rect 1800 7400 1900 7400
rect 1400 7400 1400 7400
rect 1800 7400 1800 7400
rect 1300 7400 1400 7400
rect 1700 7400 1700 7400
rect 1600 7400 1600 7400
rect 1500 7400 1600 7500
rect 1500 7500 1500 7500
rect 1500 7500 1500 7500
rect 1600 7500 1600 7500
rect 1300 7500 1300 7600
rect 1600 7500 1700 7600
rect 1400 7600 1400 7600
rect 1700 7600 1700 7600
rect 1400 7600 1500 7600
rect 1800 7600 1800 7600
rect 1500 7600 1500 7600
rect 1900 7600 1900 7600
rect 1600 7600 1600 7600
rect 1900 7600 2000 7600
rect 1700 7600 1700 7700
rect 1700 7700 1800 7700
rect 1800 7700 1800 7700
rect 1700 7700 1700 7700
rect 1600 7700 1600 7800
rect 1500 7800 1600 7800
rect 1900 7800 2000 7800
rect 1500 7800 1500 7800
rect 1900 7800 1900 7800
rect 1400 7800 1400 7800
rect 1800 7800 1800 7800
rect 1300 7800 1300 7800
rect 1700 7800 1700 7800
rect 1600 7800 1700 7900
rect 1600 7900 1600 7900
rect 1500 7900 1500 7900
rect 1400 7900 1400 7900
rect 1300 7900 1300 7900
rect 1600 8100 1700 8100
rect 1500 8100 1500 8100
rect 1800 8100 1800 8100
rect 1800 8100 1800 8100
rect 1400 8100 1400 8200
rect 1400 8200 1400 8200
rect 1900 8200 1900 8200
rect 1300 8200 1400 8200
rect 1500 8200 1600 8200
rect 1700 8200 1700 8200
rect 1400 8200 1500 8200
rect 1800 8200 1800 8200
rect 1900 8200 2000 8200
rect 1400 8200 1400 8300
rect 2000 8300 2000 8300
rect 1900 8300 1900 8300
rect 1400 8300 1400 8300
rect 1300 8300 1300 8300
rect 1900 8300 1900 8300
rect 2000 8300 2000 8300
rect 2000 8300 2000 8400
rect 1300 8500 1300 8500
rect 1400 8500 1400 8500
rect 2000 8500 2000 8500
rect 2000 8500 2000 8500
rect 1900 8500 1900 8500
rect 1900 8500 1900 8600
rect 1300 8600 1300 8600
rect 1500 8600 1600 8600
rect 2000 8600 2000 8600
rect 1900 8600 1900 8600
rect 1400 8600 1400 8600
rect 1800 8600 1900 8700
rect 1900 8700 1900 8700
rect 1500 8700 1600 8700
rect 1600 8800 1700 8800
rect 1500 8800 1500 8900
rect 1800 8800 1800 8900
rect 1800 8900 1800 8900
rect 1400 8900 1400 8900
rect 1400 8900 1400 8900
rect 1900 8900 1900 8900
rect 1300 8900 1400 9000
rect 1500 8900 1600 9000
rect 1700 8900 1700 9000
rect 1400 9000 1500 9000
rect 1800 9000 1800 9000
rect 1900 9000 2000 9000
rect 1400 9000 1400 9000
rect 2000 9000 2000 9000
rect 1900 9000 1900 9100
rect 1400 9100 1400 9100
rect 1300 9100 1300 9100
rect 1900 9100 1900 9100
rect 2000 9100 2000 9100
rect 2000 9100 2000 9100
rect 1300 9200 1300 9200
rect 1400 9200 1400 9200
rect 2000 9200 2000 9300
rect 2000 9300 2000 9300
rect 1900 9300 1900 9300
rect 1900 9300 1900 9300
rect 1300 9300 1300 9300
rect 1500 9300 1600 9400
rect 2000 9300 2000 9400
rect 1900 9400 1900 9400
rect 1400 9400 1400 9400
rect 1800 9400 1900 9400
rect 1900 9400 1900 9400
rect 1500 9400 1600 9500
rect 1800 9600 1900 9700
rect 1900 9700 1900 9700
rect 1900 9700 1900 9700
rect 1800 9700 1800 9800
rect 2000 9800 2000 9800
rect 1900 9800 1900 9800
rect 2000 9800 2000 9800
rect 1300 10400 1300 10500
rect 1400 10500 1400 10500
rect 1500 10500 1500 10500
rect 1600 10500 1600 10600
rect 1300 10600 1400 10600
rect 1400 10600 1400 10600
rect 1700 10600 1700 10600
rect 1400 10600 1500 10600
rect 1700 10600 1700 10600
rect 1500 10600 1500 10600
rect 1500 10600 1600 10700
rect 1800 10600 1800 10700
rect 2200 10600 2200 10700
rect 1600 10700 1600 10700
rect 2100 10700 2100 10700
rect 1600 10700 1700 10700
rect 1900 10700 1900 10700
rect 2000 10700 2000 10700
rect 2200 10700 2200 10700
rect 1700 10700 1700 10700
rect 2000 10700 2000 10700
rect 1700 10700 1800 10700
rect 2200 10700 2200 10700
rect 2000 10800 2100 10800
rect 1700 10800 1700 10800
rect 2000 10800 2000 10800
rect 1900 10800 2000 10800
rect 1600 10800 1600 10900
rect 1900 10800 1900 10900
rect 1800 10900 1900 10900
rect 1500 10900 1500 10900
rect 1800 10900 1800 10900
rect 1700 10900 1800 10900
rect 1400 10900 1400 10900
rect 1700 10900 1700 10900
rect 1300 11000 1300 11000
rect 1600 11000 1600 11000
rect 1500 11000 1500 11000
rect 1400 11000 1400 11100
rect 1300 11100 1300 11100
rect 1600 11200 1700 11200
rect 1500 11200 1500 11200
rect 1800 11200 1800 11200
rect 1400 11300 1400 11300
rect 1900 11300 1900 11300
rect 1500 11300 1600 11300
rect 1700 11300 1700 11300
rect 1300 11300 1300 11400
rect 1500 11300 1500 11400
rect 1800 11300 1800 11400
rect 1900 11300 2000 11400
rect 1400 11400 1400 11400
rect 1800 11400 1900 11400
rect 1300 11400 1300 11500
rect 1400 11400 1400 11500
rect 1900 11400 1900 11500
rect 2000 11400 2000 11500
rect 2800 11500 2800 11500
rect 2900 11500 3000 11500
rect 2700 11500 2700 11500
rect 3000 11500 3000 11500
rect 2600 11600 2600 11600
rect 2800 11600 2800 11600
rect 2900 11600 2900 11600
rect 1300 11600 1300 11600
rect 1400 11600 1400 11600
rect 1900 11600 1900 11600
rect 2000 11600 2000 11600
rect 2700 11600 2700 11600
rect 3000 11600 3000 11600
rect 2700 11600 2700 11600
rect 3200 11600 3200 11600
rect 2500 11600 2500 11600
rect 2600 11600 2600 11600
rect 3100 11600 3100 11600
rect 3200 11600 3200 11600
rect 2500 11600 2500 11700
rect 3200 11600 3300 11700
rect 3300 11700 3300 11700
rect 1300 11700 1300 11700
rect 1900 11700 2000 11700
rect 1600 11700 1600 11700
rect 1700 11700 1700 11700
rect 2400 11700 2400 11700
rect 1400 11800 1400 11800
rect 1900 11800 1900 11800
rect 2500 11800 2500 11800
rect 2800 11800 2900 11800
rect 3200 11800 3200 11800
rect 1400 11800 1500 11800
rect 1800 11800 1800 11800
rect 2400 11800 2400 11800
rect 2500 11800 2500 11800
rect 1600 11800 1700 11800
rect 2400 11800 2500 11900
rect 3300 11800 3300 11900
rect 3400 11800 3400 11900
rect 2800 11900 2800 11900
rect 2900 11900 2900 11900
rect 2600 11900 2600 11900
rect 3100 11900 3100 11900
rect 3300 11900 3300 11900
rect 2300 11900 2300 11900
rect 2400 11900 2400 11900
rect 3400 11900 3400 11900
rect 2300 11900 2300 12000
rect 2600 11900 2600 12000
rect 2700 11900 2700 12000
rect 3000 11900 3000 12000
rect 3100 11900 3100 12000
rect 3400 11900 3400 12000
rect 1300 12000 1800 12000
rect 1800 12000 1900 12000
rect 2600 12000 2600 12100
rect 3100 12000 3100 12100
rect 1900 12100 1900 12100
rect 2700 12100 2700 12100
rect 3000 12100 3000 12100
rect 2300 12100 2300 12100
rect 2600 12100 2600 12100
rect 3100 12100 3100 12100
rect 3400 12100 3400 12100
rect 1800 12100 1800 12100
rect 2300 12100 2300 12100
rect 3000 12100 3000 12100
rect 3300 12100 3300 12100
rect 1800 12100 1900 12200
rect 2400 12100 2400 12200
rect 3000 12100 3000 12200
rect 1900 12200 1900 12200
rect 2000 12200 2000 12200
rect 2800 12200 2800 12200
rect 2900 12200 2900 12200
rect 2000 12200 2000 12200
rect 2700 12200 2700 12200
rect 3000 12200 3000 12200
rect 3400 12200 3400 12200
rect 2300 12200 2400 12200
rect 3300 12200 3400 12200
rect 3200 12200 3300 12300
rect 2400 12300 2400 12300
rect 3100 12300 3100 12300
rect 3300 12300 3300 12300
rect 2000 12300 2000 12300
rect 2400 12300 2400 12300
rect 3200 12300 3200 12300
rect 2500 12300 2500 12300
rect 3000 12300 3000 12300
rect 2500 12300 2500 12400
rect 3100 12300 3100 12400
rect 2400 12400 2400 12400
rect 2500 12400 2600 12400
rect 3000 12400 3000 12400
rect 2400 12400 2500 12400
rect 2600 12400 2600 12400
rect 3100 12400 3100 12400
rect 2600 12400 2600 12400
rect 2900 12400 2900 12400
rect 1900 12400 1900 12500
rect 2500 12400 2500 12500
rect 2700 12400 2700 12500
rect 2900 12400 2900 12500
rect 3000 12400 3000 12500
rect 2800 12500 2800 12500
rect 3000 12500 3000 12500
rect 3000 12500 3000 12500
rect 2600 12500 2700 12500
rect 2900 12500 2900 12500
rect 2700 12500 2800 12600
rect 1300 12600 2000 12600
rect 3300 12700 3300 12700
rect 3400 12700 3400 12700
rect 3300 12800 3300 12800
rect 1400 12900 1400 12900
rect 1500 12900 1600 12900
rect 1400 12900 1400 12900
rect 1300 13000 1300 13000
rect 1400 13000 1400 13000
rect 1400 13000 1400 13000
rect 2500 13000 2600 13000
rect 1300 13100 1300 13100
rect 3000 13100 3000 13100
rect 2900 13100 3000 13100
rect 2900 13100 2900 13200
rect 1400 13200 1400 13200
rect 3000 13200 3000 13200
rect 2800 13200 2800 13300
rect 2900 13200 3000 13300
rect 2800 13300 2800 13300
rect 2800 13300 2800 13300
rect 2800 13400 2800 13400
rect 2600 13400 2700 13400
rect 2800 13400 2800 13400
rect 2600 13400 2600 13400
rect 2600 13500 2700 13500
rect 2600 13500 2600 13500
rect 1600 13600 1700 13700
rect 1500 13700 1500 13700
rect 1800 13700 1800 13700
rect 2500 13700 2500 13700
rect 1400 13700 1500 13700
rect 1800 13700 1800 13700
rect 1400 13700 1400 13700
rect 1900 13700 1900 13700
rect 2600 13700 2600 13700
rect 2700 13700 2700 13700
rect 1500 13800 1600 13800
rect 1700 13800 1700 13800
rect 2800 13800 2800 13800
rect 1500 13800 1500 13800
rect 1800 13800 1800 13800
rect 2500 13800 2600 13800
rect 2800 13800 2900 13800
rect 1300 13800 1300 13800
rect 1400 13800 1500 13800
rect 1800 13800 1800 13800
rect 2000 13800 2000 13800
rect 1400 13800 1400 13800
rect 1800 13800 1900 13800
rect 2600 13800 2700 13800
rect 2900 13800 3000 13800
rect 1400 13800 1400 13900
rect 1900 13800 1900 13900
rect 2700 13800 2700 13900
rect 3000 13800 3000 13900
rect 1300 13900 1300 13900
rect 2000 13900 2000 13900
rect 2800 13900 2800 13900
rect 1400 13900 1400 13900
rect 1900 13900 1900 13900
rect 3100 13900 3100 13900
rect 2900 13900 2900 13900
rect 3200 13900 3200 13900
rect 2900 13900 2900 13900
rect 3000 14000 3000 14000
rect 1300 14000 1300 14000
rect 2000 14000 2000 14000
rect 3000 14000 3000 14000
rect 1300 14000 1300 14100
rect 2000 14000 2000 14100
rect 2900 14000 2900 14100
rect 2800 14100 2900 14100
rect 3100 14100 3200 14100
rect 1800 14100 1800 14100
rect 2700 14100 2800 14100
rect 3000 14100 3100 14100
rect 1500 14100 1500 14100
rect 1700 14100 1800 14100
rect 2700 14100 2700 14100
rect 3000 14100 3000 14100
rect 2600 14200 2600 14200
rect 2900 14200 2900 14200
rect 2500 14200 2500 14200
rect 2800 14200 2800 14200
rect 2700 14200 2700 14200
rect 1000 14200 2000 14300
rect 2700 14200 2700 14300
rect 2600 14300 2600 14300
rect 2500 14300 2500 14300
rect 1600 14400 1700 14400
rect 2500 14400 2600 14400
rect 1500 14400 1500 14500
rect 1800 14400 1800 14500
rect 2600 14400 2600 14500
rect 1800 14500 1800 14500
rect 2700 14500 2700 14500
rect 2800 14500 2800 14500
rect 1400 14500 1400 14500
rect 2900 14500 2900 14500
rect 1400 14500 1400 14500
rect 1900 14500 1900 14500
rect 2500 14500 2500 14500
rect 2900 14500 3000 14500
rect 1300 14500 1400 14600
rect 1500 14500 1600 14600
rect 1700 14500 1700 14600
rect 2600 14500 2600 14600
rect 3000 14500 3000 14600
rect 2700 14600 2700 14600
rect 3100 14600 3100 14600
rect 1400 14600 1500 14600
rect 1800 14600 1800 14600
rect 1900 14600 2000 14600
rect 2800 14600 2800 14600
rect 3200 14600 3200 14600
rect 1400 14600 1400 14600
rect 2800 14600 2900 14600
rect 2000 14600 2000 14600
rect 2900 14600 2900 14600
rect 1900 14600 1900 14700
rect 3000 14600 3000 14700
rect 1400 14700 1400 14700
rect 3000 14700 3000 14700
rect 1300 14700 1300 14700
rect 1900 14700 1900 14700
rect 2000 14700 2000 14700
rect 2900 14700 2900 14700
rect 2000 14700 2000 14700
rect 2900 14700 2900 14700
rect 2800 14700 2800 14700
rect 3100 14700 3100 14700
rect 2700 14700 2700 14800
rect 3000 14700 3100 14800
rect 2600 14800 2600 14800
rect 3000 14800 3000 14800
rect 2500 14800 2600 14800
rect 2900 14800 2900 14800
rect 2800 14800 2800 14800
rect 1300 14800 1300 14800
rect 1400 14800 1400 14800
rect 2700 14800 2800 14800
rect 2000 14800 2000 14900
rect 2700 14800 2700 14900
rect 2000 14900 2000 14900
rect 1900 14900 1900 14900
rect 2700 14900 2700 14900
rect 1900 14900 1900 14900
rect 2800 14900 2800 14900
rect 1300 14900 1300 14900
rect 2500 14900 2500 14900
rect 2800 14900 2900 14900
rect 1500 14900 1600 15000
rect 2000 14900 2000 15000
rect 2600 14900 2600 15000
rect 2900 14900 2900 15000
rect 1900 15000 1900 15000
rect 2600 15000 2700 15000
rect 3000 15000 3000 15000
rect 1400 15000 1400 15000
rect 2700 15000 2700 15000
rect 3100 15000 3100 15000
rect 1800 15000 1900 15000
rect 2800 15000 2800 15000
rect 3100 15000 3200 15000
rect 1900 15000 1900 15000
rect 2900 15000 2900 15000
rect 1500 15000 1600 15100
rect 2900 15000 3000 15100
rect 3000 15100 3000 15100
rect 2900 15100 2900 15100
rect 2800 15100 2800 15100
rect 2700 15100 2800 15200
rect 3100 15100 3200 15200
rect 2700 15200 2700 15200
rect 3100 15200 3100 15200
rect 1800 15200 2000 15200
rect 2600 15200 2600 15200
rect 3000 15200 3000 15200
rect 1400 15200 1400 15200
rect 2500 15200 2500 15200
rect 2900 15200 2900 15200
rect 1400 15200 1400 15200
rect 1600 15200 1600 15200
rect 2000 15200 2000 15200
rect 2800 15200 2900 15200
rect 1600 15200 1600 15300
rect 1900 15200 1900 15300
rect 2800 15200 2800 15300
rect 1300 15300 1300 15300
rect 2700 15300 2700 15300
rect 2600 15300 2600 15300
rect 1300 15300 1300 15300
rect 1400 15300 1400 15300
rect 1900 15300 1900 15300
rect 2500 15300 2500 15300
rect 1400 15300 1400 15300
rect 1900 15300 1900 15300
rect 2000 15300 2000 15300
rect 1500 15300 1600 15400
rect 2000 15300 2000 15400
rect 1300 15400 1300 15400
rect 1400 15400 1400 15400
rect 1700 15400 1700 15400
rect 1600 15400 1600 15400
rect 1700 15500 1700 15500
rect 1600 15500 1600 15500
rect 1900 15500 1900 15500
rect 2000 15500 2000 15500
rect 1300 15500 1300 15500
rect 1700 15500 1700 15500
rect 1300 15500 1300 15600
rect 1600 15500 1600 15600
rect 2300 15600 2700 15600
rect 3000 15600 3200 15600
rect 1400 15600 1400 15600
rect 1800 15600 1800 15600
rect 1800 15600 1800 15600
rect 1300 15600 1300 15600
rect 1400 15600 1400 15700
rect 1600 16200 1700 16200
rect 1500 16200 1500 16200
rect 1800 16200 1800 16200
rect 1900 16200 1900 16300
rect 1300 16300 1400 16300
rect 1900 16300 1900 16300
rect 2200 16300 2200 16300
rect 1500 16300 1600 16300
rect 1700 16300 1700 16300
rect 2200 16300 2200 16300
rect 1300 16300 1300 16300
rect 1400 16300 1500 16300
rect 1800 16300 1800 16300
rect 1900 16300 2000 16300
rect 2100 16300 2100 16400
rect 1400 16400 1400 16400
rect 1800 16400 1900 16400
rect 1300 16400 1300 16400
rect 2000 16400 2000 16400
rect 2200 16400 2200 16400
rect 1400 16400 1400 16400
rect 1900 16400 1900 16400
rect 1300 16500 1300 16500
rect 2000 16500 2000 16500
rect 2100 16500 2100 16500
rect 2200 16500 2200 16500
rect 2200 16500 2200 16600
rect 1300 16600 1300 16600
rect 1900 16600 2000 16600
rect 2200 16600 2200 16600
rect 1500 16600 1500 16600
rect 1800 16600 1800 16600
rect 1500 16600 1500 16700
rect 1700 16600 1800 16700
rect 2000 16600 2000 16700
rect 2200 16600 2200 16700
rect 2100 16700 2100 16700
rect 2000 16700 2100 16800
rect 1300 16800 2000 16800
rect 1400 17100 1400 17100
rect 1500 17100 1500 17100
rect 1400 17100 1400 17100
rect 1500 17100 1500 17100
rect 1300 17100 1400 17200
rect 1300 17200 1300 17200
rect 1300 17200 1300 17200
rect 1400 17200 1400 17200
rect 1300 17300 1300 17300
rect 1400 17400 1400 17400
rect 1300 17400 1300 17400
rect 1400 17400 1500 17400
rect 1500 17400 2000 17500
rect 1400 17500 1400 17500
rect 1400 17500 1400 17500
rect 1500 17500 1500 17600
rect 1800 18200 1900 18200
rect 1900 18200 1900 18200
rect 1900 18200 1900 18200
rect 1800 18300 1800 18300
rect 2000 18300 2000 18300
rect 1900 18300 1900 18300
rect 2000 18300 2000 18300
rect 1600 18600 1700 18600
rect 1500 18600 1500 18600
rect 1800 18600 1800 18600
rect 1400 18700 1400 18700
rect 1900 18700 1900 18700
rect 1500 18700 1600 18700
rect 1700 18700 1700 18700
rect 1300 18700 1300 18800
rect 1500 18700 1500 18800
rect 1800 18700 1800 18800
rect 1900 18700 2000 18800
rect 1400 18800 1400 18800
rect 1800 18800 1900 18800
rect 1300 18800 1300 18900
rect 1400 18800 1400 18900
rect 1900 18800 1900 18900
rect 2000 18800 2000 18900
rect 1300 19000 1300 19000
rect 1400 19000 1400 19000
rect 1900 19000 1900 19000
rect 2000 19000 2000 19000
rect 1300 19100 1300 19100
rect 1900 19100 2000 19100
rect 1600 19100 1600 19100
rect 1700 19100 1700 19100
rect 1400 19200 1400 19200
rect 1900 19200 1900 19200
rect 1400 19200 1500 19200
rect 1800 19200 1800 19200
rect 1600 19200 1700 19200
rect 2500 19700 3500 19800
rect 2500 19800 3500 19800
rect 2500 19800 3500 19800
rect 2500 19800 3500 19800
rect 2500 19800 3500 19800
rect 2500 19800 3500 19900
rect 2500 19900 3500 19900
rect 2500 19900 3500 19900
rect 2500 19900 3500 19900
rect 2500 19900 3500 19900
rect 2500 19900 3500 20000
rect 2500 20000 3500 20000
rect 2500 20000 3500 20000
rect 2500 20000 3500 20000
rect 2500 20000 3500 20000
rect 2500 20000 3500 20100
rect 2500 20100 3500 20100
rect 2500 20100 3400 20100
rect 2500 20100 3400 20100
rect 2500 20100 3400 20100
rect 2500 20100 3400 20200
rect 2500 20200 3400 20200
rect 2500 20200 3400 20200
rect 2500 20200 3400 20200
rect 2500 20200 3400 20200
rect 2500 20200 3400 20300
rect 2500 20300 3400 20300
rect 2500 20300 3400 20300
rect 2500 20300 3400 20300
rect 2400 20300 3400 20300
rect 2400 20300 3400 20400
rect 2400 20400 3400 20400
rect 2400 20400 3400 20400
rect 2400 20400 3400 20400
rect 2400 20400 3400 20400
rect 2400 20400 3400 20500
rect 2400 20500 3400 20500
rect 2400 20500 3400 20500
rect 2400 20500 3400 20500
rect 2400 20500 3400 20500
rect 2400 20500 3400 20600
rect 2400 20600 3400 20600
rect 2400 20600 3400 20600
rect 2400 20600 3400 20600
rect 2400 20600 3400 20600
rect 2400 20600 3300 20700
rect 2400 20700 3300 20700
rect 2300 20700 3300 20700
rect 2300 20700 3300 20700
rect 2300 20700 3300 20700
rect 2300 20700 3300 20800
rect 2300 20800 3300 20800
rect 2300 20800 3300 20800
rect 2300 20800 3300 20800
rect 2300 20800 3300 20800
rect 2300 20800 3300 20900
rect 2300 20900 3300 20900
rect 2200 20900 3300 20900
rect 2200 20900 3300 20900
rect 2200 20900 3300 20900
rect 2200 20900 3300 21000
rect 2200 21000 3200 21000
rect 2200 21000 3200 21000
rect 2200 21000 3200 21000
rect 2200 21000 3200 21000
rect 2200 21000 3200 21100
rect 2200 21100 3200 21100
rect 2100 21100 3200 21100
rect 2100 21100 3200 21100
rect 2100 21100 3200 21100
rect 2100 21100 3200 21200
rect 2100 21200 3200 21200
rect 2100 21200 3200 21200
rect 2100 21200 3100 21200
rect 2000 21200 3100 21200
rect 2000 21200 3100 21300
rect 2000 21300 3100 21300
rect 2000 21300 3100 21300
rect 2000 21300 3100 21300
rect 2000 21300 3100 21300
rect 2000 21300 3100 21400
rect 1900 21400 3100 21400
rect 1900 21400 3100 21400
rect 1900 21400 3100 21400
rect 1900 21400 3000 21400
rect 1900 21400 3000 21500
rect 1900 21500 3000 21500
rect 1800 21500 3000 21500
rect 1800 21500 3000 21500
rect 1800 21500 3000 21500
rect 1800 21500 3000 21600
rect 1800 21600 3000 21600
rect 1700 21600 2900 21600
rect 1700 21600 2900 21600
rect 1700 21600 2900 21600
rect 1700 21600 2900 21700
rect 1700 21700 2900 21700
rect 1600 21700 2900 21700
rect 1600 21700 2900 21700
rect 1600 21700 2900 21700
rect 1500 21700 2800 21800
rect 1500 21800 2800 21800
rect 1500 21800 2800 21800
rect 1500 21800 2800 21800
rect 1500 21800 2800 21800
rect 1400 21800 2800 21900
rect 1400 21900 2800 21900
rect 1400 21900 2700 21900
rect 1300 21900 2700 21900
rect 1300 21900 2700 21900
rect 1300 21900 2700 22000
<< metal2 >>
rect 1300 7000 1300 7100
rect 1400 7100 1400 7100
rect 1500 7100 1500 7100
rect 1600 7100 1600 7100
rect 1600 7100 1700 7100
rect 1300 7100 1400 7200
rect 1700 7100 1700 7200
rect 1400 7200 1400 7200
rect 1500 7200 1500 7200
rect 1900 7200 1900 7200
rect 1600 7200 1600 7200
rect 1900 7200 2000 7200
rect 1700 7200 1700 7300
rect 1800 7300 1800 7300
rect 1800 7300 1800 7300
rect 1700 7300 1800 7300
rect 1600 7300 1600 7400
rect 1900 7300 1900 7400
rect 1500 7400 1500 7400
rect 1400 7400 1500 7400
rect 1800 7400 1800 7400
rect 1400 7400 1400 7400
rect 1700 7400 1700 7400
rect 1600 7400 1600 7400
rect 1500 7400 1500 7500
rect 1400 7500 1400 7500
rect 1500 7500 1600 7500
rect 1600 7500 1600 7600
rect 1400 7600 1400 7600
rect 1700 7600 1700 7600
rect 1500 7600 1500 7600
rect 1800 7600 1800 7600
rect 1500 7600 1600 7600
rect 1600 7600 1600 7600
rect 1900 7600 1900 7600
rect 1800 7700 1800 7700
rect 1800 7700 1800 7700
rect 1800 7700 1800 7700
rect 1700 7700 1700 7700
rect 1600 7700 1600 7800
rect 1600 7800 1600 7800
rect 1900 7800 1900 7800
rect 1500 7800 1500 7800
rect 1800 7800 1900 7800
rect 1400 7800 1400 7800
rect 1800 7800 1800 7800
rect 1300 7800 1300 7800
rect 1600 7800 1600 7900
rect 1500 7900 1600 7900
rect 1500 7900 1500 7900
rect 1400 7900 1400 7900
rect 1300 7900 1300 7900
rect 1500 8100 1500 8100
rect 1500 8100 1500 8100
rect 1800 8100 1800 8100
rect 1400 8100 1400 8100
rect 1800 8100 1900 8100
rect 1500 8200 1500 8200
rect 1700 8200 1700 8200
rect 1500 8200 1500 8200
rect 1800 8200 1800 8200
rect 1300 8200 1300 8200
rect 1300 8300 1300 8300
rect 1400 8300 1400 8300
rect 1300 8300 1300 8400
rect 1300 8400 1300 8400
rect 2000 8400 2000 8400
rect 2000 8400 2000 8400
rect 1300 8400 1300 8400
rect 1300 8400 1300 8500
rect 2000 8400 2000 8500
rect 2000 8500 2000 8500
rect 1400 8500 1400 8500
rect 1300 8500 1300 8500
rect 1500 8600 1500 8600
rect 2000 8600 2000 8600
rect 1300 8600 1400 8600
rect 1500 8600 1500 8600
rect 1400 8600 1400 8600
rect 1900 8600 2000 8600
rect 1400 8600 1400 8700
rect 1500 8700 1500 8700
rect 1600 8700 1700 8700
rect 1500 8800 1500 8900
rect 1500 8900 1500 8900
rect 1800 8900 1800 8900
rect 1400 8900 1400 8900
rect 1800 8900 1900 8900
rect 1500 8900 1500 9000
rect 1700 8900 1700 9000
rect 1500 9000 1500 9000
rect 1800 9000 1800 9000
rect 1300 9000 1300 9000
rect 1300 9000 1300 9000
rect 1400 9000 1400 9000
rect 1300 9100 1300 9100
rect 1300 9100 1300 9100
rect 2000 9100 2000 9100
rect 2000 9100 2000 9200
rect 1300 9200 1300 9200
rect 1300 9200 1300 9200
rect 2000 9200 2000 9200
rect 2000 9200 2000 9200
rect 1400 9200 1400 9300
rect 1300 9300 1300 9300
rect 1500 9300 1500 9300
rect 2000 9300 2000 9300
rect 1300 9300 1400 9400
rect 1500 9300 1500 9400
rect 1400 9400 1400 9400
rect 1900 9400 2000 9400
rect 1400 9400 1400 9400
rect 1500 9400 1500 9400
rect 1600 9400 1700 9500
rect 1800 9600 1800 9700
rect 1900 9700 2000 9700
rect 1800 9700 1800 9800
rect 1900 9800 1900 9800
rect 2000 9800 2000 9800
rect 2000 9800 2000 9800
rect 1300 10000 1400 10000
rect 1900 10000 2000 10000
rect 1300 10400 1300 10500
rect 1400 10500 1400 10500
rect 1500 10500 1500 10500
rect 1300 10500 1300 10600
rect 1500 10500 1600 10600
rect 1600 10600 1600 10600
rect 1400 10600 1400 10600
rect 1600 10600 1700 10600
rect 2200 10600 2200 10600
rect 1500 10600 1500 10600
rect 1700 10600 1800 10600
rect 2100 10600 2100 10600
rect 2200 10600 2200 10600
rect 2100 10600 2100 10700
rect 1600 10700 1600 10700
rect 1800 10700 1900 10700
rect 1900 10700 1900 10700
rect 1700 10700 1700 10700
rect 1900 10700 2000 10700
rect 2000 10700 2000 10700
rect 2200 10700 2200 10700
rect 1800 10700 1800 10800
rect 2100 10700 2100 10800
rect 1800 10800 1800 10800
rect 2100 10800 2100 10800
rect 1800 10800 1800 10800
rect 1700 10800 1800 10800
rect 2000 10800 2000 10800
rect 1700 10800 1700 10800
rect 1600 10800 1700 10900
rect 1900 10800 1900 10900
rect 1600 10900 1600 10900
rect 1800 10900 1800 10900
rect 1500 10900 1500 10900
rect 1700 10900 1700 10900
rect 1400 10900 1400 11000
rect 1600 10900 1700 11000
rect 1600 11000 1600 11000
rect 1500 11000 1600 11000
rect 1500 11000 1500 11000
rect 1400 11000 1500 11000
rect 1400 11000 1400 11100
rect 1300 11100 1400 11100
rect 1500 11200 1500 11200
rect 1800 11200 1800 11200
rect 1400 11200 1500 11300
rect 1800 11200 1800 11300
rect 1400 11300 1400 11300
rect 1900 11300 1900 11300
rect 1400 11300 1400 11300
rect 1900 11300 1900 11300
rect 1300 11300 1400 11300
rect 1500 11300 1500 11300
rect 1700 11300 1800 11300
rect 1900 11300 1900 11300
rect 1400 11400 1500 11400
rect 1800 11400 1800 11400
rect 1300 11400 1300 11400
rect 2000 11400 2000 11400
rect 1400 11400 1400 11400
rect 1900 11400 1900 11400
rect 1300 11500 1300 11500
rect 2000 11500 2000 11500
rect 1300 11500 1300 11500
rect 2000 11500 2000 11500
rect 2800 11500 2900 11500
rect 2700 11500 2700 11500
rect 3000 11500 3000 11500
rect 2600 11500 2700 11500
rect 3100 11500 3100 11500
rect 1300 11500 1300 11600
rect 2000 11500 2000 11600
rect 2600 11500 2600 11600
rect 3100 11500 3100 11600
rect 1300 11600 1300 11600
rect 2000 11600 2000 11600
rect 2800 11600 2800 11600
rect 2900 11600 3000 11600
rect 3100 11600 3200 11600
rect 2500 11600 2600 11600
rect 2600 11600 2700 11600
rect 3100 11600 3100 11600
rect 1400 11600 1400 11600
rect 1900 11600 1900 11600
rect 1300 11600 1300 11700
rect 1400 11600 1400 11700
rect 1800 11600 1900 11700
rect 2000 11600 2000 11700
rect 2600 11600 2600 11700
rect 3100 11600 3100 11700
rect 1400 11700 1500 11700
rect 1800 11700 1800 11700
rect 2600 11700 2600 11700
rect 3100 11700 3200 11700
rect 1500 11700 1500 11700
rect 1800 11700 1800 11700
rect 2500 11700 2600 11700
rect 3200 11700 3200 11700
rect 1300 11700 1400 11700
rect 1500 11700 1600 11700
rect 1700 11700 1700 11700
rect 1900 11700 1900 11700
rect 2400 11700 2400 11700
rect 2500 11700 2500 11700
rect 3200 11700 3200 11700
rect 3300 11700 3300 11700
rect 1400 11700 1400 11700
rect 1900 11700 1900 11700
rect 3200 11700 3200 11700
rect 3300 11700 3300 11700
rect 1400 11700 1400 11800
rect 1900 11700 1900 11800
rect 2400 11800 2400 11800
rect 3300 11800 3300 11800
rect 2700 11800 2800 11800
rect 3000 11800 3000 11800
rect 3200 11800 3300 11800
rect 1500 11800 1500 11800
rect 1800 11800 1800 11800
rect 2700 11800 2700 11800
rect 3000 11800 3000 11800
rect 3300 11800 3400 11800
rect 3300 11800 3300 11800
rect 2300 11900 2400 11900
rect 2600 11900 2700 11900
rect 3400 11900 3400 11900
rect 2700 11900 2800 11900
rect 3000 11900 3000 11900
rect 3300 11900 3300 11900
rect 2400 11900 2400 11900
rect 2700 11900 2700 11900
rect 3000 11900 3000 11900
rect 2300 12000 2300 12000
rect 2600 12000 2600 12000
rect 3100 12000 3100 12000
rect 3400 12000 3400 12000
rect 2300 12000 2300 12000
rect 2600 12000 2600 12000
rect 3100 12000 3100 12000
rect 3400 12000 3400 12000
rect 2300 12000 2300 12000
rect 3400 12000 3400 12000
rect 2600 12000 2600 12000
rect 3100 12000 3100 12000
rect 1900 12000 1900 12100
rect 2300 12000 2300 12100
rect 3400 12000 3400 12100
rect 2300 12100 2300 12100
rect 3400 12100 3400 12100
rect 2300 12100 2300 12100
rect 3400 12100 3400 12100
rect 1300 12100 1800 12100
rect 3000 12100 3000 12100
rect 1800 12100 1800 12100
rect 2000 12100 2000 12100
rect 2600 12100 2700 12100
rect 2700 12100 2700 12100
rect 3100 12100 3100 12100
rect 2700 12100 2700 12200
rect 2700 12100 2800 12200
rect 3000 12100 3100 12200
rect 3300 12100 3300 12200
rect 2400 12200 2400 12200
rect 2700 12200 2700 12200
rect 2800 12200 2800 12200
rect 2900 12200 3000 12200
rect 3000 12200 3000 12200
rect 3400 12200 3400 12200
rect 1900 12200 1900 12200
rect 2300 12200 2400 12200
rect 2800 12200 2900 12200
rect 2000 12200 2000 12200
rect 3100 12200 3100 12200
rect 3300 12200 3300 12200
rect 2000 12200 2000 12200
rect 2400 12200 2500 12200
rect 3100 12200 3100 12200
rect 2400 12200 2400 12300
rect 3100 12200 3100 12300
rect 2000 12300 2000 12300
rect 2500 12300 2500 12300
rect 2600 12300 3000 12300
rect 2000 12300 2000 12300
rect 2400 12300 2400 12300
rect 3200 12300 3200 12300
rect 2500 12300 2500 12300
rect 2400 12300 2400 12300
rect 3100 12300 3100 12300
rect 3300 12300 3300 12300
rect 1900 12300 1900 12400
rect 2000 12300 2000 12400
rect 3300 12300 3300 12400
rect 1900 12400 1900 12400
rect 1900 12400 2000 12400
rect 1800 12400 1900 12400
rect 1900 12400 1900 12400
rect 2500 12400 2500 12400
rect 2600 12400 2600 12400
rect 1800 12400 1800 12400
rect 1900 12400 1900 12400
rect 2500 12400 2500 12400
rect 1800 12400 1800 12500
rect 1300 12500 1700 12500
rect 1900 12500 2000 12500
rect 2700 12500 2800 12500
rect 2800 12500 2800 12500
rect 2600 12500 2600 12500
rect 2600 12500 2600 12500
rect 2900 12500 3000 12500
rect 2700 12500 2700 12500
rect 2900 12500 2900 12500
rect 3400 12600 3400 12700
rect 3400 12700 3400 12700
rect 3400 12700 3400 12700
rect 3300 12700 3300 12700
rect 3400 12700 3400 12800
rect 3300 12800 3400 12800
rect 3300 12800 3300 12800
rect 1500 12900 1500 12900
rect 1500 12900 1500 12900
rect 1300 12900 1400 13000
rect 1300 13000 1300 13000
rect 1400 13000 1400 13000
rect 3100 13000 3100 13000
rect 3000 13000 3100 13100
rect 3000 13100 3000 13100
rect 1300 13100 1300 13100
rect 1300 13100 1300 13100
rect 2900 13200 2900 13200
rect 3000 13200 3000 13200
rect 2900 13200 2900 13200
rect 3000 13200 3000 13200
rect 2900 13200 2900 13200
rect 3000 13200 3000 13200
rect 2700 13300 2800 13300
rect 2900 13300 2900 13300
rect 2700 13300 2700 13300
rect 2800 13300 2900 13300
rect 2700 13300 2700 13400
rect 2800 13300 2800 13400
rect 2600 13400 2600 13400
rect 2700 13400 2700 13500
rect 2700 13500 2700 13500
rect 2700 13500 2700 13500
rect 2500 13500 2600 13600
rect 3100 13500 3200 13600
rect 1500 13700 1500 13700
rect 1800 13700 1800 13700
rect 2500 13700 2500 13700
rect 2600 13700 2600 13700
rect 1400 13700 1400 13700
rect 1900 13700 1900 13700
rect 2700 13700 2700 13700
rect 2700 13700 2700 13800
rect 1500 13800 1500 13800
rect 1700 13800 1800 13800
rect 2500 13800 2500 13800
rect 1300 13800 1300 13800
rect 1500 13800 1500 13800
rect 1800 13800 1800 13800
rect 1900 13800 2000 13800
rect 2800 13800 2800 13800
rect 2600 13800 2600 13800
rect 2900 13800 2900 13800
rect 2700 13800 2700 13800
rect 2700 13800 2700 13900
rect 3000 13800 3000 13900
rect 1400 13900 1400 13900
rect 1900 13900 1900 13900
rect 3000 13900 3100 13900
rect 1300 13900 1300 13900
rect 2000 13900 2000 13900
rect 2800 13900 2800 13900
rect 1300 13900 1300 13900
rect 2000 13900 2000 13900
rect 2900 13900 2900 13900
rect 3100 13900 3200 13900
rect 1300 13900 1300 14000
rect 2000 13900 2000 14000
rect 3000 13900 3000 14000
rect 1300 14000 1300 14000
rect 2000 14000 2000 14000
rect 3000 14000 3100 14000
rect 3100 14000 3100 14000
rect 3000 14000 3000 14000
rect 1400 14000 1400 14000
rect 1900 14000 1900 14000
rect 3000 14000 3000 14000
rect 1300 14100 1300 14100
rect 1900 14100 2000 14100
rect 2900 14100 2900 14100
rect 2800 14100 2800 14100
rect 3100 14100 3100 14100
rect 1400 14100 1400 14100
rect 1500 14100 1500 14100
rect 1900 14100 1900 14100
rect 3000 14100 3000 14100
rect 1400 14100 1400 14100
rect 1500 14100 1500 14100
rect 1800 14100 1800 14100
rect 1900 14100 1900 14100
rect 2700 14100 2700 14100
rect 1000 14100 1400 14200
rect 1600 14100 1700 14200
rect 1900 14100 2000 14200
rect 2600 14100 2700 14200
rect 2900 14100 2900 14200
rect 2900 14200 2900 14200
rect 2500 14200 2600 14200
rect 2800 14200 2800 14200
rect 2700 14200 2700 14200
rect 2600 14300 2600 14300
rect 2500 14300 2600 14300
rect 2500 14400 2500 14400
rect 1500 14400 1500 14500
rect 2600 14400 2600 14500
rect 1500 14500 1500 14500
rect 1800 14500 1800 14500
rect 2700 14500 2700 14500
rect 1400 14500 1400 14500
rect 1800 14500 1900 14500
rect 2800 14500 2800 14500
rect 2800 14500 2900 14500
rect 2500 14500 2600 14500
rect 2900 14500 2900 14500
rect 1500 14500 1500 14600
rect 1700 14500 1700 14600
rect 2600 14500 2600 14600
rect 1500 14600 1500 14600
rect 1800 14600 1800 14600
rect 2700 14600 2700 14600
rect 3100 14600 3100 14600
rect 1300 14600 1300 14600
rect 2800 14600 2800 14600
rect 3100 14600 3200 14600
rect 1300 14600 1300 14600
rect 1400 14600 1400 14600
rect 2900 14600 2900 14600
rect 3000 14600 3000 14700
rect 3000 14700 3000 14700
rect 2900 14700 3000 14700
rect 1300 14700 1300 14700
rect 1300 14700 1300 14700
rect 2000 14700 2000 14700
rect 2800 14700 2800 14700
rect 3100 14700 3100 14700
rect 2000 14700 2000 14800
rect 2700 14700 2700 14800
rect 2600 14800 2700 14800
rect 3000 14800 3000 14800
rect 1300 14800 1300 14800
rect 2600 14800 2600 14800
rect 2900 14800 2900 14800
rect 1300 14800 1300 14800
rect 2000 14800 2000 14800
rect 2800 14800 2800 14800
rect 2000 14800 2000 14800
rect 2700 14800 2700 14800
rect 1400 14800 1400 14900
rect 2600 14900 2600 14900
rect 1300 14900 1300 14900
rect 2700 14900 2800 14900
rect 1500 14900 1500 14900
rect 2000 14900 2000 14900
rect 2800 14900 2800 14900
rect 1300 14900 1400 15000
rect 1500 14900 1500 15000
rect 2600 14900 2600 15000
rect 2900 14900 2900 15000
rect 1400 15000 1400 15000
rect 2700 15000 2700 15000
rect 3000 15000 3000 15000
rect 1900 15000 2000 15000
rect 2700 15000 2800 15000
rect 1400 15000 1400 15000
rect 2800 15000 2800 15000
rect 3100 15000 3100 15000
rect 1500 15000 1500 15000
rect 1600 15000 1700 15100
rect 3000 15000 3000 15100
rect 3000 15100 3000 15100
rect 3000 15100 3000 15100
rect 2900 15100 2900 15100
rect 2800 15100 2800 15100
rect 2800 15100 2800 15200
rect 3100 15100 3100 15200
rect 2700 15200 2700 15200
rect 3000 15200 3100 15200
rect 2600 15200 2600 15200
rect 3000 15200 3000 15200
rect 1500 15200 1600 15200
rect 2500 15200 2500 15200
rect 2800 15200 2800 15200
rect 1300 15200 1400 15300
rect 2000 15200 2000 15300
rect 2700 15200 2800 15300
rect 2700 15300 2700 15300
rect 1600 15300 1600 15300
rect 2600 15300 2600 15300
rect 1500 15300 1500 15300
rect 2500 15300 2500 15300
rect 1500 15300 1600 15300
rect 1600 15300 1700 15300
rect 1400 15300 1400 15400
rect 2000 15400 2000 15400
rect 1300 15400 1300 15400
rect 1600 15400 1600 15400
rect 2000 15400 2000 15400
rect 1300 15400 1300 15400
rect 1700 15400 1700 15400
rect 2000 15400 2000 15400
rect 1300 15400 1300 15400
rect 2000 15400 2000 15500
rect 1300 15500 1300 15500
rect 1600 15500 1600 15500
rect 2000 15500 2000 15500
rect 1300 15500 1300 15500
rect 1700 15500 1700 15500
rect 2000 15500 2000 15500
rect 1300 15500 1300 15500
rect 1900 15500 1900 15500
rect 1700 15600 1700 15600
rect 2000 15600 2000 15600
rect 1600 15600 1600 15600
rect 1700 15600 1800 15600
rect 1400 15600 1400 15600
rect 1900 15600 2000 15600
rect 1600 15600 1700 15600
rect 1700 15600 1700 15700
rect 1700 15700 1700 15700
rect 1900 15700 1900 15700
rect 2900 15700 2900 15700
rect 1700 15700 1700 15700
rect 1800 15700 1900 15700
rect 1500 16200 1500 16200
rect 1700 16200 1800 16200
rect 1400 16200 1500 16200
rect 1800 16200 1800 16200
rect 1400 16200 1400 16200
rect 1800 16200 1900 16200
rect 2100 16300 2100 16300
rect 2200 16300 2200 16300
rect 1500 16300 1500 16300
rect 1800 16300 1800 16300
rect 2200 16300 2200 16300
rect 1400 16400 1400 16400
rect 1900 16400 1900 16400
rect 1300 16400 1300 16400
rect 2000 16400 2000 16400
rect 2200 16400 2200 16400
rect 1300 16400 1300 16400
rect 2000 16400 2000 16400
rect 2200 16400 2200 16400
rect 2200 16400 2200 16500
rect 1300 16500 1300 16500
rect 2000 16500 2000 16500
rect 1300 16500 1300 16500
rect 2000 16500 2000 16500
rect 2200 16500 2200 16500
rect 2200 16500 2200 16500
rect 1400 16500 1400 16600
rect 1900 16500 1900 16600
rect 2100 16500 2100 16600
rect 1300 16600 1300 16600
rect 1400 16600 1400 16600
rect 1800 16600 1900 16600
rect 1900 16600 1900 16600
rect 2100 16600 2100 16600
rect 1400 16600 1400 16600
rect 1800 16600 1800 16600
rect 2100 16600 2100 16600
rect 1400 16600 1400 16600
rect 1900 16600 1900 16600
rect 2100 16600 2100 16600
rect 1400 16600 1400 16700
rect 1900 16600 1900 16700
rect 2000 16600 2000 16700
rect 1300 16700 1400 16700
rect 1600 16700 1700 16700
rect 1900 16700 1900 16700
rect 2200 16700 2200 16700
rect 2100 16700 2200 16700
rect 2100 16700 2100 16700
rect 2000 16700 2000 16800
rect 1500 17100 1500 17100
rect 1400 17100 1400 17200
rect 1400 17200 1400 17200
rect 1300 17300 1300 17300
rect 1300 17300 1300 17300
rect 1300 17300 1300 17400
rect 1300 17400 1300 17400
rect 1300 17400 1300 17400
rect 1500 17400 1500 17500
rect 1300 17500 1300 17500
rect 1300 17500 1400 17500
rect 1500 17500 1500 17600
rect 1800 18200 1800 18200
rect 1900 18300 2000 18300
rect 1800 18300 1800 18300
rect 1900 18300 1900 18300
rect 2000 18300 2000 18400
rect 2000 18400 2000 18400
rect 1300 18500 1400 18500
rect 1900 18500 2000 18500
rect 1500 18600 1500 18600
rect 1800 18600 1800 18600
rect 1400 18600 1500 18700
rect 1800 18600 1800 18700
rect 1400 18700 1400 18700
rect 1900 18700 1900 18700
rect 1400 18700 1400 18700
rect 1900 18700 1900 18700
rect 1300 18700 1400 18700
rect 1500 18700 1500 18700
rect 1700 18700 1800 18700
rect 1900 18700 1900 18700
rect 1400 18800 1500 18800
rect 1800 18800 1800 18800
rect 1300 18800 1300 18800
rect 2000 18800 2000 18800
rect 1400 18800 1400 18800
rect 1900 18800 1900 18800
rect 1300 18900 1300 18900
rect 2000 18900 2000 18900
rect 1300 18900 1300 18900
rect 2000 18900 2000 18900
rect 1300 18900 1300 19000
rect 2000 18900 2000 19000
rect 1300 19000 1300 19000
rect 2000 19000 2000 19000
rect 1400 19000 1400 19000
rect 1900 19000 1900 19000
rect 1300 19000 1300 19100
rect 1400 19000 1400 19100
rect 1800 19000 1900 19100
rect 2000 19000 2000 19100
rect 1400 19100 1500 19100
rect 1800 19100 1800 19100
rect 1500 19100 1500 19100
rect 1800 19100 1800 19100
rect 1300 19100 1400 19100
rect 1500 19100 1600 19100
rect 1700 19100 1700 19100
rect 1900 19100 1900 19100
rect 1400 19100 1400 19100
rect 1900 19100 1900 19100
rect 1400 19100 1400 19200
rect 1900 19100 1900 19200
rect 1500 19200 1500 19200
rect 1800 19200 1800 19200
rect 1500 19700 2500 19800
rect 1500 19800 2500 19800
rect 1500 19800 2500 19800
rect 1500 19800 2500 19800
rect 1500 19800 2500 19800
rect 1500 19800 2500 19900
rect 1500 19900 2500 19900
rect 1500 19900 2500 19900
rect 1500 19900 2500 19900
rect 1500 19900 2500 19900
rect 1500 19900 2500 20000
rect 1500 20000 2500 20000
rect 1500 20000 2500 20000
rect 1500 20000 2500 20000
rect 1500 20000 2500 20000
rect 1500 20000 2500 20100
rect 1500 20100 2500 20100
rect 1500 20100 2500 20100
rect 1500 20100 2500 20100
rect 1400 20100 2500 20100
rect 1400 20100 2500 20200
rect 1400 20200 2500 20200
rect 1400 20200 2500 20200
rect 1400 20200 2500 20200
rect 1400 20200 2500 20200
rect 1400 20200 2500 20300
rect 1400 20300 2500 20300
rect 1400 20300 2500 20300
rect 1400 20300 2500 20300
rect 1400 20300 2400 20300
rect 1400 20300 2400 20400
rect 1400 20400 2400 20400
rect 1300 20400 2400 20400
rect 1300 20400 2400 20400
rect 1300 20400 2400 20400
rect 1300 20400 2400 20500
rect 1300 20500 2400 20500
rect 1300 20500 2400 20500
rect 1300 20500 2400 20500
rect 1300 20500 2400 20500
rect 1300 20500 2400 20600
rect 1300 20600 2400 20600
rect 1200 20600 2400 20600
rect 1200 20600 2400 20600
rect 1200 20600 2400 20600
rect 1200 20600 2400 20700
rect 1200 20700 2400 20700
rect 1200 20700 2300 20700
rect 1200 20700 2300 20700
rect 1100 20700 2300 20700
rect 1100 20700 2300 20800
rect 1100 20800 2300 20800
rect 1100 20800 2300 20800
rect 1100 20800 2300 20800
rect 1000 20800 2300 20800
rect 1000 20800 2300 20900
rect 1000 20900 2300 20900
rect 1000 20900 2200 20900
rect 1000 20900 2200 20900
rect 900 20900 2200 20900
rect 900 20900 2200 21000
rect 900 21000 2200 21000
rect 900 21000 2200 21000
rect 800 21000 2200 21000
rect 800 21000 2200 21000
rect 800 21000 2200 21100
rect 700 21100 2200 21100
rect 700 21100 2100 21100
rect 700 21100 2100 21100
rect 600 21100 2100 21100
rect 600 21100 2100 21200
rect 600 21200 2100 21200
rect 500 21200 2100 21200
rect 500 21200 2100 21200
rect 400 21200 2000 21200
rect 300 21200 2000 21300
rect 200 21300 200 21300
rect 200 21300 2000 21300
rect 0 21300 0 21300
rect 100 21300 2000 21300
rect 0 21300 2000 21300
rect 0 21300 2000 21300
rect 0 21300 2000 21400
rect 0 21400 1900 21400
rect 0 21400 1900 21400
rect 0 21400 1900 21400
rect 0 21400 1900 21400
rect 0 21400 1900 21500
rect 0 21500 1900 21500
rect 0 21500 1800 21500
rect 0 21500 1800 21500
rect 0 21500 1800 21500
rect 0 21500 1800 21600
rect 0 21600 1800 21600
rect 0 21600 1700 21600
rect 0 21600 1700 21600
rect 0 21600 1700 21600
rect 0 21600 1700 21700
rect 0 21700 1700 21700
rect 0 21700 1600 21700
rect 0 21700 1600 21700
rect 0 21700 1600 21700
rect 0 21700 1500 21800
rect 0 21800 1500 21800
rect 0 21800 1500 21800
rect 0 21800 1500 21800
rect 0 21800 1500 21800
rect 0 21800 1400 21900
rect 0 21900 1400 21900
rect 0 21900 1400 21900
rect 0 21900 1300 21900
rect 0 21900 1300 21900
rect 0 21900 1300 22000
<< metal3 >>
rect 500 19700 1500 19800
rect 500 19800 1500 19800
rect 500 19800 1500 19800
rect 500 19800 1500 19800
rect 500 19800 1500 19800
rect 500 19800 1500 19900
rect 500 19900 1500 19900
rect 500 19900 1500 19900
rect 500 19900 1500 19900
rect 400 19900 1500 19900
rect 400 19900 1500 20000
rect 400 20000 1500 20000
rect 400 20000 1500 20000
rect 400 20000 1500 20000
rect 400 20000 1500 20000
rect 400 20000 1500 20100
rect 400 20100 1500 20100
rect 400 20100 1500 20100
rect 300 20100 1500 20100
rect 300 20100 1400 20100
rect 300 20100 1400 20200
rect 300 20200 1400 20200
rect 200 20200 1400 20200
rect 200 20200 1400 20200
rect 200 20200 1400 20200
rect 100 20200 1400 20300
rect 100 20300 1400 20300
rect 0 20300 1400 20300
rect 0 20300 1400 20300
rect 0 20300 1400 20300
rect 0 20300 1400 20400
rect 0 20400 1400 20400
rect 0 20400 1300 20400
rect 0 20400 1300 20400
rect 0 20400 1300 20400
rect 0 20400 1300 20500
rect 0 20500 1300 20500
rect 0 20500 1300 20500
rect 0 20500 1300 20500
rect 0 20500 1300 20500
rect 0 20500 1300 20600
rect 0 20600 1300 20600
rect 0 20600 1200 20600
rect 0 20600 1200 20600
rect 0 20600 1200 20600
rect 0 20600 1200 20700
rect 0 20700 1200 20700
rect 0 20700 1200 20700
rect 0 20700 1200 20700
rect 0 20700 1100 20700
rect 0 20700 1100 20800
rect 0 20800 1100 20800
rect 0 20800 1100 20800
rect 0 20800 1100 20800
rect 0 20800 1000 20800
rect 0 20800 1000 20900
rect 0 20900 1000 20900
rect 0 20900 1000 20900
rect 0 20900 1000 20900
rect 0 20900 900 20900
rect 0 20900 900 21000
rect 0 21000 900 21000
rect 0 21000 900 21000
rect 0 21000 800 21000
rect 0 21000 800 21000
rect 0 21000 800 21100
rect 0 21100 700 21100
rect 0 21100 700 21100
rect 0 21100 700 21100
rect 0 21100 600 21100
rect 0 21100 600 21200
rect 0 21200 600 21200
rect 0 21200 500 21200
rect 0 21200 500 21200
rect 0 21200 400 21200
rect 0 21200 300 21300
rect 0 21300 200 21300
rect 200 21300 200 21300
rect 0 21300 0 21300
rect 0 21300 100 21300
<< metal4 >>
rect 2200 800 2700 800
rect 2000 800 2000 800
rect 2000 800 2900 800
rect 1900 800 3000 800
rect 1800 800 3100 900
rect 1800 900 3100 900
rect 1700 900 3200 900
rect 1700 900 3300 900
rect 1600 900 3300 900
rect 1500 900 3400 1000
rect 1500 1000 3400 1000
rect 1500 1000 3500 1000
rect 1400 1000 3500 1000
rect 1400 1000 3500 1000
rect 1300 1000 3600 1100
rect 1300 1100 3600 1100
rect 1300 1100 3700 1100
rect 1200 1100 3700 1100
rect 1200 1100 3700 1100
rect 1200 1100 3800 1200
rect 1100 1200 3800 1200
rect 1100 1200 3800 1200
rect 1100 1200 3800 1200
rect 1000 1200 3900 1200
rect 1000 1200 3900 1300
rect 1000 1300 3900 1300
rect 1000 1300 3900 1300
rect 900 1300 4000 1300
rect 900 1300 4000 1300
rect 900 1300 4000 1400
rect 900 1400 4000 1400
rect 800 1400 4100 1400
rect 800 1400 4100 1400
rect 800 1400 4100 1400
rect 800 1400 4100 1500
rect 800 1500 4200 1500
rect 700 1500 4200 1500
rect 700 1500 4200 1500
rect 700 1500 4200 1500
rect 700 1500 4200 1600
rect 700 1600 4200 1600
rect 600 1600 4300 1600
rect 600 1600 2200 1600
rect 2700 1600 4300 1600
rect 600 1600 2100 1600
rect 2800 1600 4300 1600
rect 600 1600 2000 1700
rect 2900 1600 4300 1700
rect 600 1700 2000 1700
rect 2900 1700 4300 1700
rect 600 1700 1900 1700
rect 3000 1700 4300 1700
rect 500 1700 1900 1700
rect 3000 1700 4400 1700
rect 500 1700 1800 1700
rect 3100 1700 4400 1700
rect 500 1700 1800 1800
rect 3100 1700 4400 1800
rect 500 1800 1700 1800
rect 3200 1800 4400 1800
rect 500 1800 1700 1800
rect 3200 1800 4400 1800
rect 500 1800 1700 1800
rect 3200 1800 4400 1800
rect 500 1800 1600 1800
rect 3300 1800 4400 1800
rect 400 1800 1600 1900
rect 3300 1800 4500 1900
rect 400 1900 1600 1900
rect 3300 1900 4500 1900
rect 400 1900 1500 1900
rect 3300 1900 4500 1900
rect 400 1900 1500 1900
rect 3400 1900 4500 1900
rect 400 1900 1500 1900
rect 3400 1900 4500 1900
rect 400 1900 1500 2000
rect 3400 1900 4500 2000
rect 400 2000 1400 2000
rect 3400 2000 4500 2000
rect 400 2000 1400 2000
rect 3500 2000 4500 2000
rect 400 2000 1400 2000
rect 2400 2000 2500 2000
rect 3500 2000 4600 2000
rect 300 2000 1400 2000
rect 2200 2000 2600 2000
rect 3500 2000 4600 2000
rect 300 2000 1400 2100
rect 2200 2000 2700 2100
rect 3500 2000 4600 2100
rect 300 2100 1300 2100
rect 2100 2100 2800 2100
rect 3500 2100 4600 2100
rect 300 2100 1300 2100
rect 2000 2100 2900 2100
rect 3600 2100 4600 2100
rect 300 2100 1300 2100
rect 2000 2100 2900 2100
rect 3600 2100 4600 2100
rect 300 2100 1300 2100
rect 1900 2100 2900 2100
rect 3600 2100 4600 2100
rect 300 2100 1300 2200
rect 1900 2100 3000 2200
rect 3600 2100 4600 2200
rect 300 2200 1200 2200
rect 1900 2200 3000 2200
rect 3600 2200 4600 2200
rect 300 2200 1200 2200
rect 1800 2200 3000 2200
rect 3700 2200 4600 2200
rect 300 2200 1200 2200
rect 1800 2200 3100 2200
rect 3700 2200 4700 2200
rect 200 2200 1200 2200
rect 1800 2200 3100 2200
rect 3700 2200 4700 2200
rect 200 2200 1200 2300
rect 1800 2200 3100 2300
rect 3700 2200 4700 2300
rect 200 2300 1200 2300
rect 1700 2300 3200 2300
rect 3700 2300 4700 2300
rect 200 2300 1200 2300
rect 1700 2300 3200 2300
rect 3700 2300 4700 2300
rect 200 2300 1100 2300
rect 1700 2300 3200 2300
rect 3700 2300 4700 2300
rect 200 2300 1100 2300
rect 1700 2300 3200 2300
rect 3700 2300 4700 2300
rect 200 2300 1100 2400
rect 1600 2300 3200 2400
rect 3800 2300 4700 2400
rect 200 2400 1100 2400
rect 1600 2400 3300 2400
rect 3800 2400 4700 2400
rect 200 2400 1100 2400
rect 1600 2400 3300 2400
rect 3800 2400 4700 2400
rect 200 2400 1100 2400
rect 1600 2400 3300 2400
rect 3800 2400 4700 2400
rect 200 2400 1100 2400
rect 1600 2400 3300 2400
rect 3800 2400 4700 2400
rect 200 2400 1100 2500
rect 1600 2400 3300 2500
rect 3800 2400 4700 2500
rect 200 2500 1100 2500
rect 1500 2500 3300 2500
rect 3800 2500 4800 2500
rect 200 2500 1100 2500
rect 1500 2500 3300 2500
rect 3800 2500 4800 2500
rect 100 2500 1000 2500
rect 1500 2500 3400 2500
rect 3800 2500 4800 2500
rect 100 2500 1000 2500
rect 1500 2500 3400 2500
rect 3800 2500 4800 2500
rect 100 2500 1000 2600
rect 1500 2500 3400 2600
rect 3900 2500 4800 2600
rect 100 2600 1000 2600
rect 1500 2600 3400 2600
rect 3900 2600 4800 2600
rect 100 2600 1000 2600
rect 1500 2600 3400 2600
rect 3900 2600 4800 2600
rect 100 2600 1000 2600
rect 1500 2600 3400 2600
rect 3900 2600 4800 2600
rect 100 2600 1000 2600
rect 1400 2600 3400 2600
rect 3900 2600 4800 2600
rect 100 2600 1000 2700
rect 1400 2600 3400 2700
rect 3900 2600 4800 2700
rect 100 2700 1000 2700
rect 1400 2700 3400 2700
rect 3900 2700 4800 2700
rect 100 2700 1000 2700
rect 1400 2700 3500 2700
rect 3900 2700 4800 2700
rect 100 2700 1000 2700
rect 1400 2700 3500 2700
rect 3900 2700 4800 2700
rect 100 2700 1000 2700
rect 1400 2700 3500 2700
rect 3900 2700 4800 2700
rect 100 2700 1000 2800
rect 1400 2700 3500 2800
rect 3900 2700 4800 2800
rect 100 2800 1000 2800
rect 1400 2800 3500 2800
rect 3900 2800 4800 2800
rect 100 2800 1000 2800
rect 1400 2800 3500 2800
rect 3900 2800 4800 2800
rect 100 2800 1000 2800
rect 1400 2800 3500 2800
rect 3900 2800 4800 2800
rect 100 2800 1000 2800
rect 1400 2800 3500 2800
rect 3900 2800 4800 2800
rect 100 2800 1000 2900
rect 1400 2800 3500 2900
rect 3900 2800 4800 2900
rect 100 2900 1100 2900
rect 1400 2900 3500 2900
rect 3900 2900 4800 2900
rect 100 2900 1100 2900
rect 1400 2900 3500 2900
rect 3900 2900 4800 2900
rect 100 2900 1100 2900
rect 1400 2900 3500 2900
rect 3900 2900 4800 2900
rect 100 2900 1200 2900
rect 1300 2900 3500 2900
rect 3900 2900 4800 2900
rect 100 2900 1200 3000
rect 1300 2900 3500 3000
rect 3900 2900 4800 3000
rect 100 3000 1300 3000
rect 1300 3000 3500 3000
rect 3800 3000 4800 3000
rect 100 3000 3500 3000
rect 3800 3000 4800 3000
rect 100 3000 3500 3000
rect 3700 3000 4800 3000
rect 100 3000 3500 3000
rect 3700 3000 4900 3000
rect 100 3000 4900 3100
rect 100 3100 4900 3100
rect 100 3100 4900 3100
rect 100 3100 4900 3100
rect 100 3100 4900 3100
rect 100 3100 4900 3200
rect 100 3200 4900 3200
rect 100 3200 4900 3200
rect 100 3200 4900 3200
rect 100 3200 4900 3200
rect 100 3200 4900 3300
rect 100 3300 4900 3300
rect 100 3300 4900 3300
rect 100 3300 4900 3300
rect 100 3300 4900 3300
rect 100 3300 4800 3400
rect 100 3400 4800 3400
rect 100 3400 4800 3400
rect 100 3400 4800 3400
rect 100 3400 4800 3400
rect 100 3400 4800 3500
rect 100 3500 4800 3500
rect 100 3500 4800 3500
rect 100 3500 1500 3500
rect 1700 3500 3200 3500
rect 3400 3500 4800 3500
rect 100 3500 1400 3500
rect 1800 3500 3100 3500
rect 3500 3500 4800 3500
rect 100 3500 1400 3600
rect 1800 3500 3100 3600
rect 3500 3500 4800 3600
rect 100 3600 1300 3600
rect 1800 3600 3100 3600
rect 3600 3600 4800 3600
rect 100 3600 1300 3600
rect 1900 3600 3000 3600
rect 3600 3600 4800 3600
rect 100 3600 1300 3600
rect 1900 3600 3000 3600
rect 3600 3600 4800 3600
rect 100 3600 1300 3600
rect 1900 3600 3000 3600
rect 3600 3600 4800 3600
rect 100 3600 1300 3700
rect 1900 3600 3000 3700
rect 3700 3600 4800 3700
rect 100 3700 1200 3700
rect 1900 3700 3000 3700
rect 3700 3700 4800 3700
rect 100 3700 1200 3700
rect 2000 3700 3000 3700
rect 3700 3700 4800 3700
rect 100 3700 1200 3700
rect 2000 3700 2900 3700
rect 3700 3700 4800 3700
rect 100 3700 1200 3700
rect 2000 3700 2900 3700
rect 3700 3700 4800 3700
rect 100 3700 1200 3800
rect 2000 3700 2900 3800
rect 3700 3700 4800 3800
rect 100 3800 1200 3800
rect 2000 3800 2900 3800
rect 3700 3800 4800 3800
rect 100 3800 1200 3800
rect 2000 3800 2900 3800
rect 3700 3800 4800 3800
rect 100 3800 1200 3800
rect 2000 3800 2900 3800
rect 3700 3800 4800 3800
rect 100 3800 1200 3800
rect 2000 3800 2900 3800
rect 3700 3800 4800 3800
rect 100 3800 1200 3900
rect 2000 3800 2900 3900
rect 3700 3800 4800 3900
rect 200 3900 1200 3900
rect 2000 3900 2900 3900
rect 3800 3900 4800 3900
rect 200 3900 1200 3900
rect 2000 3900 2900 3900
rect 3800 3900 4800 3900
rect 200 3900 1200 3900
rect 2000 3900 2900 3900
rect 3800 3900 4700 3900
rect 200 3900 1200 3900
rect 2000 3900 2900 3900
rect 3800 3900 4700 3900
rect 200 3900 1200 4000
rect 2000 3900 2900 4000
rect 3800 3900 4700 4000
rect 200 4000 1200 4000
rect 2000 4000 2900 4000
rect 3800 4000 4700 4000
rect 200 4000 1200 4000
rect 2000 4000 2900 4000
rect 3700 4000 4700 4000
rect 200 4000 1200 4000
rect 2000 4000 2900 4000
rect 3700 4000 4700 4000
rect 200 4000 1200 4000
rect 2000 4000 2900 4000
rect 3700 4000 4700 4000
rect 200 4000 1200 4100
rect 2000 4000 2900 4100
rect 3700 4000 4700 4100
rect 200 4100 1200 4100
rect 2000 4100 2900 4100
rect 3700 4100 4700 4100
rect 200 4100 1200 4100
rect 2000 4100 2900 4100
rect 3700 4100 4700 4100
rect 200 4100 1200 4100
rect 2000 4100 2900 4100
rect 3700 4100 4700 4100
rect 200 4100 1200 4100
rect 2000 4100 2900 4100
rect 3700 4100 4700 4100
rect 300 4100 1200 4200
rect 2000 4100 2900 4200
rect 3700 4100 4700 4200
rect 300 4200 1200 4200
rect 1900 4200 3000 4200
rect 3700 4200 4600 4200
rect 300 4200 1200 4200
rect 1900 4200 3000 4200
rect 3700 4200 4600 4200
rect 300 4200 1300 4200
rect 1900 4200 3000 4200
rect 3600 4200 4600 4200
rect 300 4200 1300 4200
rect 1900 4200 3000 4200
rect 3600 4200 4600 4200
rect 300 4200 1300 4300
rect 1900 4200 3000 4300
rect 3600 4200 4600 4300
rect 300 4300 1300 4300
rect 1900 4300 3100 4300
rect 3600 4300 4600 4300
rect 300 4300 1400 4300
rect 1800 4300 3100 4300
rect 3600 4300 4600 4300
rect 300 4300 1400 4300
rect 1800 4300 3100 4300
rect 3500 4300 4600 4300
rect 300 4300 1400 4300
rect 1700 4300 3200 4300
rect 3500 4300 4600 4300
rect 400 4300 1500 4400
rect 1700 4300 3300 4400
rect 3400 4300 4600 4400
rect 400 4400 4500 4400
rect 400 4400 4500 4400
rect 400 4400 4500 4400
rect 400 4400 4500 4400
rect 400 4400 4500 4500
rect 400 4500 4500 4500
rect 400 4500 4500 4500
rect 500 4500 4500 4500
rect 500 4500 4400 4500
rect 500 4500 4400 4600
rect 500 4600 4400 4600
rect 500 4600 4400 4600
rect 500 4600 4400 4600
rect 500 4600 4400 4600
rect 600 4600 4400 4700
rect 600 4700 4300 4700
rect 600 4700 4300 4700
rect 600 4700 4300 4700
rect 600 4700 4300 4700
rect 600 4700 4300 4800
rect 700 4800 4300 4800
rect 700 4800 4200 4800
rect 700 4800 4200 4800
rect 700 4800 4200 4800
rect 700 4800 4200 4900
rect 700 4900 4200 4900
rect 800 4900 4100 4900
rect 800 4900 4100 4900
rect 800 4900 4100 4900
rect 800 4900 4100 5000
rect 900 5000 4100 5000
rect 900 5000 4000 5000
rect 900 5000 4000 5000
rect 900 5000 4000 5000
rect 1000 5000 4000 5100
rect 1000 5100 3900 5100
rect 1000 5100 3900 5100
rect 1000 5100 3900 5100
rect 1100 5100 3900 5100
rect 1100 5100 3800 5200
rect 1100 5200 3800 5200
rect 1100 5200 3800 5200
rect 1200 5200 3700 5200
rect 1200 5200 3700 5200
rect 1200 5200 3700 5300
rect 1300 5300 3600 5300
rect 1300 5300 3600 5300
rect 1300 5300 3600 5300
rect 1400 5300 3500 5300
rect 1400 5300 3500 5400
rect 1500 5400 3400 5400
rect 1500 5400 3400 5400
rect 1600 5400 3300 5400
rect 1600 5400 3300 5400
rect 1700 5400 3200 5500
rect 1700 5500 3200 5500
rect 1800 5500 3100 5500
rect 1900 5500 3000 5500
rect 2000 5500 3000 5500
rect 2100 5500 2100 5600
rect 2100 5500 2800 5600
rect 2300 5600 2600 5600
rect 1100 6400 1200 6400
rect 1100 6400 1200 6500
rect 1100 6500 1200 6500
rect 1100 6500 1200 6500
rect 1100 6500 1200 6500
rect 1100 6500 1200 6500
rect 1100 6500 1200 6600
rect 1100 6600 1200 6600
rect 1100 6600 1200 6600
rect 1100 6600 1200 6600
rect 1100 6600 1200 6600
rect 1100 6600 1200 6700
rect 1100 6700 1200 6700
rect 1100 6700 1200 6700
rect 1100 6700 1200 6700
rect 1100 6700 1200 6700
rect 1100 6700 2000 6800
rect 1100 6800 2000 6800
rect 1100 6800 2000 6800
rect 1100 6800 2000 6800
rect 1100 6800 2000 6800
rect 1100 6800 2000 6900
rect 1100 6900 1200 6900
rect 1100 6900 1200 6900
rect 1100 6900 1200 6900
rect 1100 6900 1200 6900
rect 1100 6900 1200 7000
rect 1100 7000 1200 7000
rect 1100 7000 1200 7000
rect 1100 7000 1200 7000
rect 1100 7000 1200 7000
rect 1100 7000 1200 7100
rect 1300 7000 1300 7100
rect 1100 7100 1200 7100
rect 1300 7100 1400 7100
rect 1100 7100 1200 7100
rect 1300 7100 1500 7100
rect 1100 7100 1200 7100
rect 1300 7100 1600 7100
rect 1100 7100 1200 7100
rect 1300 7100 1600 7100
rect 1100 7100 1200 7200
rect 1400 7100 1700 7200
rect 1100 7200 1200 7200
rect 1400 7200 1800 7200
rect 1500 7200 1900 7200
rect 1600 7200 1900 7200
rect 1700 7200 2000 7200
rect 1700 7200 2000 7300
rect 1800 7300 2000 7300
rect 1800 7300 2000 7300
rect 1800 7300 2000 7300
rect 1700 7300 2000 7300
rect 1600 7300 1900 7400
rect 1500 7400 1800 7400
rect 1500 7400 1800 7400
rect 1400 7400 1700 7400
rect 1300 7400 1600 7400
rect 1300 7400 1500 7500
rect 1300 7500 1500 7500
rect 1300 7500 1400 7500
rect 1300 7500 1500 7500
rect 1300 7500 1500 7500
rect 1300 7500 1600 7600
rect 1400 7600 1700 7600
rect 1500 7600 1800 7600
rect 1600 7600 1900 7600
rect 1600 7600 1900 7600
rect 1700 7600 2000 7700
rect 1800 7700 2000 7700
rect 1800 7700 2000 7700
rect 1800 7700 2000 7700
rect 1700 7700 2000 7700
rect 1600 7700 2000 7800
rect 1600 7800 1900 7800
rect 1500 7800 1800 7800
rect 1400 7800 1800 7800
rect 1300 7800 1700 7800
rect 1300 7800 1600 7900
rect 1300 7900 1500 7900
rect 1300 7900 1500 7900
rect 1300 7900 1400 7900
rect 1500 8100 1800 8100
rect 1500 8100 1800 8100
rect 1400 8100 1800 8100
rect 1400 8100 1900 8200
rect 1400 8200 1900 8200
rect 1400 8200 1500 8200
rect 1600 8200 1700 8200
rect 1700 8200 1900 8200
rect 1300 8200 1500 8200
rect 1600 8200 1700 8200
rect 1800 8200 1900 8200
rect 1300 8200 1400 8200
rect 1600 8200 1700 8200
rect 1800 8200 1900 8200
rect 1300 8200 1400 8300
rect 1600 8200 1700 8300
rect 1800 8200 2000 8300
rect 1300 8300 1400 8300
rect 1600 8300 1700 8300
rect 1900 8300 2000 8300
rect 1300 8300 1400 8300
rect 1600 8300 1700 8300
rect 1900 8300 2000 8300
rect 1300 8300 1400 8300
rect 1600 8300 1700 8300
rect 1900 8300 2000 8300
rect 1300 8300 1400 8300
rect 1600 8300 1700 8300
rect 1900 8300 2000 8300
rect 1300 8300 1400 8400
rect 1600 8300 1700 8400
rect 1900 8300 2000 8400
rect 1300 8400 1400 8400
rect 1600 8400 1700 8400
rect 1900 8400 2000 8400
rect 1300 8400 1400 8400
rect 1600 8400 1700 8400
rect 1900 8400 2000 8400
rect 1300 8400 1400 8400
rect 1600 8400 1700 8400
rect 1900 8400 2000 8400
rect 1300 8400 1400 8400
rect 1600 8400 1700 8400
rect 1900 8400 2000 8400
rect 1300 8400 1400 8500
rect 1600 8400 1700 8500
rect 1900 8400 2000 8500
rect 1300 8500 1400 8500
rect 1600 8500 1700 8500
rect 1900 8500 2000 8500
rect 1300 8500 1400 8500
rect 1600 8500 1700 8500
rect 1900 8500 2000 8500
rect 1300 8500 1400 8500
rect 1600 8500 1700 8500
rect 1900 8500 2000 8500
rect 1300 8500 1400 8500
rect 1600 8500 1700 8500
rect 1900 8500 2000 8500
rect 1300 8500 1400 8600
rect 1600 8500 1700 8600
rect 1900 8500 2000 8600
rect 1300 8600 1500 8600
rect 1600 8600 1700 8600
rect 1900 8600 2000 8600
rect 1400 8600 1500 8600
rect 1600 8600 1700 8600
rect 1900 8600 2000 8600
rect 1400 8600 1700 8600
rect 1900 8600 2000 8600
rect 1400 8600 1700 8600
rect 1900 8600 1900 8600
rect 1400 8600 1700 8700
rect 1900 8600 1900 8700
rect 1500 8700 1700 8700
rect 1500 8800 1800 8900
rect 1500 8900 1800 8900
rect 1400 8900 1800 8900
rect 1400 8900 1900 8900
rect 1400 8900 1900 8900
rect 1400 8900 1500 9000
rect 1600 8900 1700 9000
rect 1700 8900 1900 9000
rect 1300 9000 1500 9000
rect 1600 9000 1700 9000
rect 1800 9000 1900 9000
rect 1300 9000 1400 9000
rect 1600 9000 1700 9000
rect 1800 9000 1900 9000
rect 1300 9000 1400 9000
rect 1600 9000 1700 9000
rect 1800 9000 2000 9000
rect 1300 9000 1400 9000
rect 1600 9000 1700 9000
rect 1900 9000 2000 9000
rect 1300 9000 1400 9100
rect 1600 9000 1700 9100
rect 1900 9000 2000 9100
rect 1300 9100 1400 9100
rect 1600 9100 1700 9100
rect 1900 9100 2000 9100
rect 1300 9100 1400 9100
rect 1600 9100 1700 9100
rect 1900 9100 2000 9100
rect 1300 9100 1400 9100
rect 1600 9100 1700 9100
rect 1900 9100 2000 9100
rect 1300 9100 1400 9100
rect 1600 9100 1700 9100
rect 1900 9100 2000 9100
rect 1300 9100 1400 9200
rect 1600 9100 1700 9200
rect 1900 9100 2000 9200
rect 1300 9200 1400 9200
rect 1600 9200 1700 9200
rect 1900 9200 2000 9200
rect 1300 9200 1400 9200
rect 1600 9200 1700 9200
rect 1900 9200 2000 9200
rect 1300 9200 1400 9200
rect 1600 9200 1700 9200
rect 1900 9200 2000 9200
rect 1300 9200 1400 9200
rect 1600 9200 1700 9200
rect 1900 9200 2000 9200
rect 1300 9200 1400 9300
rect 1600 9200 1700 9300
rect 1900 9200 2000 9300
rect 1300 9300 1400 9300
rect 1600 9300 1700 9300
rect 1900 9300 2000 9300
rect 1300 9300 1400 9300
rect 1600 9300 1700 9300
rect 1900 9300 2000 9300
rect 1300 9300 1400 9300
rect 1600 9300 1700 9300
rect 1900 9300 2000 9300
rect 1300 9300 1500 9300
rect 1600 9300 1700 9300
rect 1900 9300 2000 9300
rect 1400 9300 1500 9400
rect 1600 9300 1700 9400
rect 1900 9300 2000 9400
rect 1400 9400 1700 9400
rect 1900 9400 2000 9400
rect 1400 9400 1700 9400
rect 1900 9400 1900 9400
rect 1400 9400 1700 9400
rect 1900 9400 1900 9400
rect 1500 9400 1700 9400
rect 1300 9600 1400 9600
rect 1300 9600 1400 9600
rect 1300 9600 1400 9600
rect 1300 9600 1400 9600
rect 1100 9600 1800 9700
rect 1100 9700 1900 9700
rect 1100 9700 1900 9700
rect 1100 9700 1900 9700
rect 1100 9700 1900 9700
rect 1300 9700 1400 9800
rect 1800 9700 2000 9800
rect 1300 9800 1400 9800
rect 1900 9800 2000 9800
rect 1300 9800 1400 9800
rect 1900 9800 2000 9800
rect 1300 9800 1400 9800
rect 1900 9800 2000 9800
rect 1300 9800 1400 9800
rect 1900 9800 2000 9800
rect 1300 9800 1400 9900
rect 1900 9800 2000 9900
rect 1300 9900 1400 9900
rect 1900 9900 2000 9900
rect 1300 9900 1400 9900
rect 1900 9900 2000 9900
rect 1300 9900 1400 9900
rect 1900 9900 2000 9900
rect 1300 9900 1400 9900
rect 1900 9900 2000 9900
rect 1300 9900 1400 10000
rect 1900 9900 2000 10000
rect 1300 10500 1400 10500
rect 1300 10500 1400 10500
rect 1300 10500 1500 10500
rect 2100 10500 2200 10500
rect 1300 10500 1500 10500
rect 2100 10500 2200 10500
rect 1300 10500 1500 10600
rect 2100 10500 2200 10600
rect 1400 10600 1600 10600
rect 2100 10600 2200 10600
rect 1400 10600 1600 10600
rect 2100 10600 2200 10600
rect 1500 10600 1700 10600
rect 2100 10600 2200 10600
rect 1500 10600 1700 10600
rect 2100 10600 2200 10600
rect 1600 10600 1800 10700
rect 2100 10600 2200 10700
rect 1600 10700 1800 10700
rect 2100 10700 2200 10700
rect 1700 10700 1900 10700
rect 2000 10700 2200 10700
rect 1700 10700 1900 10700
rect 2000 10700 2200 10700
rect 1800 10700 2200 10700
rect 1800 10700 2100 10800
rect 1800 10800 2100 10800
rect 1800 10800 2000 10800
rect 1800 10800 2000 10800
rect 1700 10800 1900 10800
rect 1700 10800 1900 10900
rect 1600 10900 1800 10900
rect 1500 10900 1800 10900
rect 1500 10900 1700 10900
rect 1400 10900 1700 10900
rect 1400 10900 1600 11000
rect 1300 11000 1600 11000
rect 1300 11000 1500 11000
rect 1300 11000 1500 11000
rect 1300 11000 1400 11000
rect 1300 11000 1400 11100
rect 1300 11100 1300 11100
rect 1500 11200 1800 11200
rect 1500 11200 1800 11300
rect 1400 11300 1900 11300
rect 1400 11300 1900 11300
rect 1400 11300 1900 11300
rect 1400 11300 1500 11300
rect 1800 11300 1900 11300
rect 1300 11300 1500 11400
rect 1800 11300 1900 11400
rect 1300 11400 1400 11400
rect 1800 11400 2000 11400
rect 1300 11400 1400 11400
rect 1900 11400 2000 11400
rect 1300 11400 1400 11400
rect 1900 11400 2000 11400
rect 1300 11400 1400 11400
rect 1900 11400 2000 11400
rect 1300 11400 1400 11500
rect 1900 11400 2000 11500
rect 1300 11500 1400 11500
rect 1900 11500 2000 11500
rect 1300 11500 1400 11500
rect 1900 11500 2000 11500
rect 1300 11500 1400 11500
rect 1900 11500 2000 11500
rect 2700 11500 3000 11500
rect 1300 11500 1400 11500
rect 1900 11500 2000 11500
rect 2700 11500 3100 11500
rect 1300 11500 1400 11600
rect 1900 11500 2000 11600
rect 2600 11500 3100 11600
rect 1300 11600 1400 11600
rect 1900 11600 2000 11600
rect 2600 11600 2800 11600
rect 3000 11600 3100 11600
rect 1300 11600 1400 11600
rect 1900 11600 2000 11600
rect 2600 11600 2700 11600
rect 3000 11600 3200 11600
rect 1300 11600 1400 11600
rect 1900 11600 2000 11600
rect 2500 11600 2600 11600
rect 3100 11600 3200 11600
rect 1300 11600 1400 11600
rect 1900 11600 2000 11600
rect 2500 11600 2600 11600
rect 3100 11600 3200 11600
rect 1300 11600 1400 11700
rect 1900 11600 2000 11700
rect 2500 11600 2600 11700
rect 3100 11600 3200 11700
rect 1300 11700 1400 11700
rect 1800 11700 2000 11700
rect 2500 11700 2600 11700
rect 3200 11700 3300 11700
rect 1300 11700 1500 11700
rect 1800 11700 1900 11700
rect 2400 11700 2500 11700
rect 3200 11700 3300 11700
rect 1400 11700 1500 11700
rect 1700 11700 1900 11700
rect 2400 11700 2500 11700
rect 3200 11700 3300 11700
rect 1400 11700 1900 11700
rect 2400 11700 2500 11700
rect 3200 11700 3300 11700
rect 1400 11700 1900 11800
rect 2400 11700 2500 11800
rect 3200 11700 3300 11800
rect 1400 11800 1900 11800
rect 2400 11800 2500 11800
rect 3200 11800 3300 11800
rect 1500 11800 1800 11800
rect 2400 11800 2500 11800
rect 2800 11800 3000 11800
rect 3300 11800 3300 11800
rect 1500 11800 1800 11800
rect 2400 11800 2500 11800
rect 2700 11800 3000 11800
rect 3300 11800 3300 11800
rect 2400 11800 2500 11800
rect 2700 11800 3000 11800
rect 3300 11800 3400 11800
rect 2400 11800 2400 11900
rect 2700 11800 3100 11900
rect 3300 11800 3400 11900
rect 2400 11900 2400 11900
rect 2700 11900 2800 11900
rect 2900 11900 3100 11900
rect 3300 11900 3400 11900
rect 2300 11900 2400 11900
rect 2600 11900 2700 11900
rect 3000 11900 3100 11900
rect 3300 11900 3400 11900
rect 2300 11900 2400 11900
rect 2600 11900 2700 11900
rect 3000 11900 3100 11900
rect 3300 11900 3400 11900
rect 2300 11900 2400 11900
rect 2600 11900 2700 11900
rect 3000 11900 3100 11900
rect 3300 11900 3400 11900
rect 2300 11900 2400 12000
rect 2600 11900 2700 12000
rect 3000 11900 3100 12000
rect 3300 11900 3400 12000
rect 2300 12000 2400 12000
rect 2600 12000 2700 12000
rect 3000 12000 3100 12000
rect 3300 12000 3400 12000
rect 2300 12000 2400 12000
rect 2600 12000 2700 12000
rect 3000 12000 3100 12000
rect 3300 12000 3400 12000
rect 2300 12000 2400 12000
rect 2600 12000 2700 12000
rect 3000 12000 3100 12000
rect 3300 12000 3400 12000
rect 1300 12000 1800 12000
rect 2300 12000 2400 12000
rect 2600 12000 2700 12000
rect 3000 12000 3100 12000
rect 3300 12000 3400 12000
rect 1300 12000 1900 12100
rect 2300 12000 2400 12100
rect 2600 12000 2700 12100
rect 3000 12000 3100 12100
rect 3300 12000 3400 12100
rect 1300 12100 1900 12100
rect 2300 12100 2400 12100
rect 2600 12100 2700 12100
rect 3000 12100 3100 12100
rect 3300 12100 3400 12100
rect 1300 12100 1900 12100
rect 2300 12100 2400 12100
rect 2600 12100 2700 12100
rect 3000 12100 3100 12100
rect 3300 12100 3400 12100
rect 1800 12100 2000 12100
rect 2300 12100 2400 12100
rect 2600 12100 2700 12100
rect 3000 12100 3100 12100
rect 3300 12100 3400 12100
rect 1800 12100 2000 12100
rect 2300 12100 2400 12100
rect 2700 12100 2700 12100
rect 3000 12100 3100 12100
rect 3300 12100 3400 12100
rect 1900 12100 2000 12200
rect 2300 12100 2400 12200
rect 2700 12100 2700 12200
rect 3000 12100 3000 12200
rect 3300 12100 3400 12200
rect 1900 12200 2000 12200
rect 2300 12200 2400 12200
rect 2700 12200 2800 12200
rect 3000 12200 3000 12200
rect 3300 12200 3400 12200
rect 1900 12200 2000 12200
rect 2400 12200 2400 12200
rect 2700 12200 2800 12200
rect 2900 12200 3000 12200
rect 3300 12200 3400 12200
rect 1900 12200 2000 12200
rect 2400 12200 2400 12200
rect 2600 12200 3100 12200
rect 3300 12200 3400 12200
rect 1900 12200 2000 12200
rect 2400 12200 2400 12200
rect 2600 12200 3100 12200
rect 3300 12200 3300 12200
rect 1900 12200 2000 12300
rect 2400 12200 2500 12300
rect 2600 12200 3100 12300
rect 3300 12200 3300 12300
rect 1900 12300 2000 12300
rect 2400 12300 2500 12300
rect 3000 12300 3100 12300
rect 3200 12300 3300 12300
rect 1900 12300 2000 12300
rect 2400 12300 2500 12300
rect 3000 12300 3100 12300
rect 3200 12300 3300 12300
rect 1900 12300 2000 12300
rect 2400 12300 2500 12300
rect 3000 12300 3100 12300
rect 3200 12300 3300 12300
rect 1900 12300 2000 12300
rect 2400 12300 2500 12300
rect 3000 12300 3100 12300
rect 3200 12300 3300 12300
rect 1900 12300 2000 12400
rect 2400 12300 2500 12400
rect 3000 12300 3100 12400
rect 3200 12300 3300 12400
rect 1900 12400 2000 12400
rect 2400 12400 2500 12400
rect 3000 12400 3100 12400
rect 1900 12400 1900 12400
rect 2500 12400 2600 12400
rect 3000 12400 3100 12400
rect 1900 12400 1900 12400
rect 2500 12400 2600 12400
rect 3000 12400 3100 12400
rect 1800 12400 1900 12400
rect 2500 12400 2600 12400
rect 2900 12400 3000 12400
rect 1800 12400 1900 12500
rect 2500 12400 2700 12500
rect 2900 12400 3000 12500
rect 1700 12500 1900 12500
rect 2500 12500 2700 12500
rect 2800 12500 3000 12500
rect 1300 12500 2000 12500
rect 2600 12500 3000 12500
rect 1300 12500 2000 12500
rect 2600 12500 2900 12500
rect 1300 12500 2000 12500
rect 2700 12500 2900 12500
rect 1300 12500 2000 12600
rect 3300 12600 3400 12600
rect 3300 12600 3400 12600
rect 3300 12600 3400 12700
rect 3300 12700 3400 12700
rect 3300 12700 3400 12700
rect 3300 12700 3400 12700
rect 3300 12700 3400 12700
rect 2200 12700 2400 12800
rect 2500 12700 3400 12800
rect 2200 12800 2400 12800
rect 2500 12800 3400 12800
rect 2200 12800 2400 12800
rect 2500 12800 3400 12800
rect 1300 12800 2000 12800
rect 2200 12800 2400 12800
rect 2500 12800 3300 12800
rect 1300 12800 2000 12800
rect 2200 12800 2400 12800
rect 2500 12800 3300 12800
rect 1300 12800 2000 12900
rect 1300 12900 2000 12900
rect 1300 12900 2000 12900
rect 1400 12900 1500 12900
rect 1400 12900 1500 12900
rect 1400 12900 1400 13000
rect 1300 13000 1400 13000
rect 1300 13000 1400 13000
rect 1300 13000 1400 13000
rect 1300 13000 1400 13000
rect 3100 13000 3200 13000
rect 1300 13000 1400 13100
rect 2500 13000 2600 13100
rect 3100 13000 3200 13100
rect 1300 13100 1400 13100
rect 2500 13100 2600 13100
rect 3000 13100 3200 13100
rect 1300 13100 1400 13100
rect 2500 13100 2600 13100
rect 3000 13100 3200 13100
rect 1300 13100 1400 13100
rect 2500 13100 2600 13100
rect 3000 13100 3200 13100
rect 1300 13100 1400 13100
rect 2500 13100 2600 13100
rect 3000 13100 3200 13100
rect 1300 13100 1400 13200
rect 2500 13100 2600 13200
rect 2900 13100 3100 13200
rect 3100 13100 3200 13200
rect 1300 13200 1400 13200
rect 2500 13200 2600 13200
rect 2900 13200 3000 13200
rect 3100 13200 3200 13200
rect 2500 13200 2600 13200
rect 2900 13200 3000 13200
rect 3100 13200 3200 13200
rect 2500 13200 2600 13200
rect 2900 13200 3000 13200
rect 3100 13200 3200 13200
rect 2500 13200 2600 13200
rect 2800 13200 3000 13200
rect 3100 13200 3200 13200
rect 2500 13200 2600 13300
rect 2800 13200 2900 13300
rect 3100 13200 3200 13300
rect 2500 13300 2600 13300
rect 2800 13300 2900 13300
rect 3100 13300 3200 13300
rect 2500 13300 2600 13300
rect 2800 13300 2900 13300
rect 3100 13300 3200 13300
rect 2500 13300 2600 13300
rect 2800 13300 2900 13300
rect 3100 13300 3200 13300
rect 2500 13300 2600 13300
rect 2700 13300 2800 13300
rect 3100 13300 3200 13300
rect 2500 13300 2600 13400
rect 2700 13300 2800 13400
rect 3100 13300 3200 13400
rect 2500 13400 2600 13400
rect 2700 13400 2800 13400
rect 3100 13400 3200 13400
rect 2500 13400 2600 13400
rect 2700 13400 2800 13400
rect 3100 13400 3200 13400
rect 2500 13400 2600 13400
rect 2600 13400 2800 13400
rect 3100 13400 3200 13400
rect 2500 13400 2600 13400
rect 2600 13400 2700 13400
rect 3100 13400 3200 13400
rect 2500 13400 2700 13500
rect 3100 13400 3200 13500
rect 2500 13500 2700 13500
rect 3100 13500 3200 13500
rect 2500 13500 2700 13500
rect 3100 13500 3200 13500
rect 2500 13500 2600 13500
rect 3100 13500 3200 13500
rect 2500 13500 2600 13500
rect 3100 13500 3200 13500
rect 1500 13700 1800 13700
rect 1500 13700 1800 13700
rect 2500 13700 2600 13700
rect 1400 13700 1900 13700
rect 2500 13700 2600 13700
rect 1400 13700 1900 13700
rect 2500 13700 2700 13700
rect 1400 13700 1900 13800
rect 2500 13700 2700 13800
rect 1300 13800 1500 13800
rect 1800 13800 1900 13800
rect 2500 13800 2800 13800
rect 1300 13800 1500 13800
rect 1800 13800 1900 13800
rect 2600 13800 2800 13800
rect 1300 13800 1400 13800
rect 1800 13800 2000 13800
rect 2600 13800 2900 13800
rect 1300 13800 1400 13800
rect 1900 13800 2000 13800
rect 2700 13800 2900 13800
rect 1300 13800 1400 13900
rect 1900 13800 2000 13900
rect 2700 13800 3000 13900
rect 1300 13900 1400 13900
rect 1900 13900 2000 13900
rect 2800 13900 3000 13900
rect 1300 13900 1400 13900
rect 1900 13900 2000 13900
rect 2800 13900 3100 13900
rect 1300 13900 1400 13900
rect 1900 13900 2000 13900
rect 2900 13900 3100 13900
rect 1300 13900 1400 13900
rect 1900 13900 2000 13900
rect 2900 13900 3200 13900
rect 1300 13900 1400 14000
rect 1900 13900 2000 14000
rect 3000 13900 3200 14000
rect 1300 14000 1400 14000
rect 1900 14000 2000 14000
rect 3100 14000 3200 14000
rect 1300 14000 1400 14000
rect 1900 14000 2000 14000
rect 3100 14000 3200 14000
rect 1300 14000 1400 14000
rect 1900 14000 2000 14000
rect 3000 14000 3200 14000
rect 1300 14000 1400 14000
rect 1900 14000 2000 14000
rect 3000 14000 3200 14000
rect 1300 14000 1400 14100
rect 1900 14000 2000 14100
rect 2900 14000 3200 14100
rect 1300 14100 1400 14100
rect 1900 14100 1900 14100
rect 2900 14100 3100 14100
rect 1300 14100 1400 14100
rect 1800 14100 1900 14100
rect 2800 14100 3100 14100
rect 1400 14100 1500 14100
rect 1800 14100 1900 14100
rect 2800 14100 3000 14100
rect 1400 14100 1500 14100
rect 1800 14100 1900 14100
rect 2700 14100 3000 14100
rect 1400 14100 1600 14200
rect 1700 14100 1900 14200
rect 2700 14100 2900 14200
rect 1000 14200 2000 14200
rect 2600 14200 2900 14200
rect 1000 14200 2000 14200
rect 2600 14200 2800 14200
rect 1000 14200 2000 14200
rect 2500 14200 2800 14200
rect 1000 14200 2000 14200
rect 2500 14200 2700 14200
rect 2500 14200 2700 14300
rect 2500 14300 2600 14300
rect 2500 14300 2500 14300
rect 2500 14400 2500 14400
rect 1500 14400 1800 14500
rect 2500 14400 2600 14500
rect 1500 14500 1800 14500
rect 2500 14500 2700 14500
rect 1400 14500 1800 14500
rect 2500 14500 2800 14500
rect 1400 14500 1900 14500
rect 2500 14500 2800 14500
rect 1400 14500 1900 14500
rect 2600 14500 2900 14500
rect 1400 14500 1500 14600
rect 1600 14500 1700 14600
rect 1700 14500 1900 14600
rect 2600 14500 3000 14600
rect 1300 14600 1500 14600
rect 1600 14600 1700 14600
rect 1800 14600 1900 14600
rect 2700 14600 3100 14600
rect 1300 14600 1400 14600
rect 1600 14600 1700 14600
rect 1800 14600 1900 14600
rect 2800 14600 3100 14600
rect 1300 14600 1400 14600
rect 1600 14600 1700 14600
rect 1800 14600 2000 14600
rect 2900 14600 3200 14600
rect 1300 14600 1400 14600
rect 1600 14600 1700 14600
rect 1900 14600 2000 14600
rect 2900 14600 3200 14600
rect 1300 14600 1400 14700
rect 1600 14600 1700 14700
rect 1900 14600 2000 14700
rect 3000 14600 3200 14700
rect 1300 14700 1400 14700
rect 1600 14700 1700 14700
rect 1900 14700 2000 14700
rect 3000 14700 3200 14700
rect 1300 14700 1400 14700
rect 1600 14700 1700 14700
rect 1900 14700 2000 14700
rect 3000 14700 3200 14700
rect 1300 14700 1400 14700
rect 1600 14700 1700 14700
rect 1900 14700 2000 14700
rect 2900 14700 3200 14700
rect 1300 14700 1400 14700
rect 1600 14700 1700 14700
rect 1900 14700 2000 14700
rect 2800 14700 3100 14700
rect 1300 14700 1400 14800
rect 1600 14700 1700 14800
rect 1900 14700 2000 14800
rect 2700 14700 3000 14800
rect 1300 14800 1400 14800
rect 1600 14800 1700 14800
rect 1900 14800 2000 14800
rect 2700 14800 3000 14800
rect 1300 14800 1400 14800
rect 1600 14800 1700 14800
rect 1900 14800 2000 14800
rect 2600 14800 2900 14800
rect 1300 14800 1400 14800
rect 1600 14800 1700 14800
rect 1900 14800 2000 14800
rect 2500 14800 2800 14800
rect 1300 14800 1400 14800
rect 1600 14800 1700 14800
rect 1900 14800 2000 14800
rect 2500 14800 2700 14800
rect 1300 14800 1400 14900
rect 1600 14800 1700 14900
rect 1900 14800 2000 14900
rect 2500 14800 2700 14900
rect 1300 14900 1400 14900
rect 1600 14900 1700 14900
rect 1900 14900 2000 14900
rect 2500 14900 2600 14900
rect 1300 14900 1400 14900
rect 1600 14900 1700 14900
rect 1900 14900 2000 14900
rect 2500 14900 2700 14900
rect 1300 14900 1400 14900
rect 1600 14900 1700 14900
rect 1900 14900 2000 14900
rect 2500 14900 2700 14900
rect 1300 14900 1500 14900
rect 1600 14900 1700 14900
rect 1900 14900 2000 14900
rect 2500 14900 2800 14900
rect 1400 14900 1500 15000
rect 1600 14900 1700 15000
rect 1900 14900 2000 15000
rect 2600 14900 2900 15000
rect 1400 15000 1700 15000
rect 1900 15000 2000 15000
rect 2700 15000 3000 15000
rect 1400 15000 1700 15000
rect 1900 15000 1900 15000
rect 2800 15000 3100 15000
rect 1400 15000 1700 15000
rect 1900 15000 1900 15000
rect 2800 15000 3100 15000
rect 1500 15000 1700 15000
rect 2900 15000 3200 15000
rect 3000 15000 3200 15100
rect 3000 15100 3200 15100
rect 3000 15100 3200 15100
rect 2900 15100 3200 15100
rect 2800 15100 3200 15100
rect 2800 15100 3100 15200
rect 2700 15200 3000 15200
rect 2600 15200 3000 15200
rect 1400 15200 1500 15200
rect 1900 15200 2000 15200
rect 2500 15200 2900 15200
rect 1400 15200 1600 15200
rect 1900 15200 2000 15200
rect 2500 15200 2800 15200
rect 1400 15200 1600 15300
rect 1900 15200 2000 15300
rect 2500 15200 2700 15300
rect 1300 15300 1600 15300
rect 1900 15300 2000 15300
rect 2500 15300 2700 15300
rect 1300 15300 1600 15300
rect 1900 15300 2000 15300
rect 2500 15300 2600 15300
rect 1300 15300 1400 15300
rect 1500 15300 1600 15300
rect 1900 15300 2000 15300
rect 1300 15300 1400 15300
rect 1600 15300 1600 15300
rect 1900 15300 2000 15300
rect 1300 15300 1400 15400
rect 1600 15300 1700 15400
rect 1900 15300 2000 15400
rect 1300 15400 1400 15400
rect 1600 15400 1700 15400
rect 1900 15400 2000 15400
rect 1300 15400 1400 15400
rect 1600 15400 1700 15400
rect 1900 15400 2000 15400
rect 1300 15400 1400 15400
rect 1600 15400 1700 15400
rect 1900 15400 2000 15400
rect 1300 15400 1400 15400
rect 1600 15400 1700 15400
rect 1900 15400 2000 15400
rect 1300 15400 1400 15500
rect 1600 15400 1700 15500
rect 1900 15400 2000 15500
rect 1300 15500 1400 15500
rect 1600 15500 1700 15500
rect 1900 15500 2000 15500
rect 1300 15500 1400 15500
rect 1600 15500 1700 15500
rect 1900 15500 2000 15500
rect 1300 15500 1400 15500
rect 1600 15500 1700 15500
rect 1900 15500 2000 15500
rect 1300 15500 1400 15500
rect 1600 15500 1700 15500
rect 1900 15500 2000 15500
rect 1300 15500 1400 15600
rect 1600 15500 1700 15600
rect 1900 15500 2000 15600
rect 1300 15600 1400 15600
rect 1600 15600 1700 15600
rect 1900 15600 2000 15600
rect 1300 15600 1400 15600
rect 1600 15600 1700 15600
rect 1800 15600 2000 15600
rect 2300 15600 2900 15600
rect 3000 15600 3200 15600
rect 1300 15600 1400 15600
rect 1600 15600 1900 15600
rect 2300 15600 2900 15600
rect 3000 15600 3200 15600
rect 1300 15600 1400 15600
rect 1700 15600 1900 15600
rect 2300 15600 2900 15600
rect 3000 15600 3200 15600
rect 1300 15600 1400 15700
rect 1700 15600 1900 15700
rect 2300 15600 2900 15700
rect 3000 15600 3200 15700
rect 1700 15700 1900 15700
rect 2300 15700 2900 15700
rect 3000 15700 3200 15700
rect 1700 15700 1800 15700
rect 1000 15900 1200 15900
rect 1300 15900 2000 15900
rect 1000 15900 1200 15900
rect 1300 15900 2000 15900
rect 1000 15900 1200 15900
rect 1300 15900 2000 15900
rect 1000 15900 1200 16000
rect 1300 15900 2000 16000
rect 1000 16000 1200 16000
rect 1300 16000 2000 16000
rect 1500 16200 1700 16200
rect 1500 16200 1800 16200
rect 1400 16200 1800 16200
rect 1400 16200 1900 16300
rect 1400 16300 1900 16300
rect 2100 16300 2200 16300
rect 1300 16300 1500 16300
rect 1700 16300 1900 16300
rect 2100 16300 2200 16300
rect 1300 16300 1500 16300
rect 1800 16300 1900 16300
rect 2100 16300 2200 16300
rect 1300 16300 1400 16300
rect 1800 16300 1900 16300
rect 2100 16300 2200 16300
rect 1300 16300 1400 16400
rect 1800 16300 2000 16400
rect 2100 16300 2200 16400
rect 1300 16400 1400 16400
rect 1900 16400 2000 16400
rect 2100 16400 2200 16400
rect 1300 16400 1400 16400
rect 1900 16400 2000 16400
rect 2100 16400 2200 16400
rect 1300 16400 1400 16400
rect 1900 16400 2000 16400
rect 2100 16400 2200 16400
rect 1300 16400 1400 16400
rect 1900 16400 2000 16400
rect 2100 16400 2200 16400
rect 1300 16400 1400 16500
rect 1900 16400 2000 16500
rect 2100 16400 2200 16500
rect 1300 16500 1400 16500
rect 1900 16500 2000 16500
rect 2100 16500 2200 16500
rect 1300 16500 1400 16500
rect 1900 16500 2000 16500
rect 2100 16500 2200 16500
rect 1300 16500 1400 16500
rect 1900 16500 2000 16500
rect 2100 16500 2200 16500
rect 1300 16500 1400 16500
rect 1900 16500 2000 16500
rect 2100 16500 2200 16500
rect 1300 16500 1400 16600
rect 1900 16500 2000 16600
rect 2100 16500 2200 16600
rect 1300 16600 1400 16600
rect 1900 16600 1900 16600
rect 2100 16600 2200 16600
rect 1300 16600 1400 16600
rect 1900 16600 1900 16600
rect 2100 16600 2200 16600
rect 1300 16600 1400 16600
rect 1800 16600 1900 16600
rect 2100 16600 2200 16600
rect 1400 16600 1500 16600
rect 1800 16600 1900 16600
rect 2100 16600 2200 16600
rect 1400 16600 1500 16700
rect 1800 16600 1900 16700
rect 2000 16600 2200 16700
rect 1400 16700 1600 16700
rect 1700 16700 1900 16700
rect 1900 16700 2200 16700
rect 1300 16700 2100 16700
rect 1300 16700 2100 16700
rect 1300 16700 2100 16700
rect 1300 16700 2000 16800
rect 1300 17000 2000 17000
rect 1300 17000 2000 17000
rect 1300 17000 2000 17100
rect 1300 17100 2000 17100
rect 1300 17100 2000 17100
rect 1400 17100 1500 17100
rect 1400 17100 1500 17100
rect 1400 17100 1400 17200
rect 1300 17200 1400 17200
rect 1300 17200 1400 17200
rect 1300 17200 1400 17200
rect 1300 17200 1400 17200
rect 1300 17200 1400 17300
rect 1300 17300 1400 17300
rect 1300 17300 1400 17300
rect 1300 17300 1400 17300
rect 1300 17300 1400 17300
rect 1300 17300 1400 17400
rect 1300 17400 1400 17400
rect 1300 17400 1400 17400
rect 1300 17400 1400 17400
rect 1300 17400 1400 17400
rect 1300 17400 1500 17500
rect 1300 17500 2000 17500
rect 1400 17500 2000 17500
rect 1400 17500 2000 17500
rect 1400 17500 2000 17500
rect 1500 17500 2000 17600
rect 1300 18100 1400 18100
rect 1300 18100 1400 18100
rect 1300 18100 1400 18200
rect 1300 18200 1400 18200
rect 1100 18200 1800 18200
rect 1100 18200 1900 18200
rect 1100 18200 1900 18200
rect 1100 18200 1900 18300
rect 1100 18300 1900 18300
rect 1300 18300 1400 18300
rect 1800 18300 2000 18300
rect 1300 18300 1400 18300
rect 1900 18300 2000 18300
rect 1300 18300 1400 18300
rect 1900 18300 2000 18300
rect 1300 18300 1400 18400
rect 1900 18300 2000 18400
rect 1300 18400 1400 18400
rect 1900 18400 2000 18400
rect 1300 18400 1400 18400
rect 1900 18400 2000 18400
rect 1300 18400 1400 18400
rect 1900 18400 2000 18400
rect 1300 18400 1400 18400
rect 1900 18400 2000 18400
rect 1300 18400 1400 18500
rect 1900 18400 2000 18500
rect 1300 18500 1400 18500
rect 1900 18500 2000 18500
rect 1300 18500 1400 18500
rect 1900 18500 2000 18500
rect 1500 18600 1800 18600
rect 1500 18600 1800 18700
rect 1400 18700 1900 18700
rect 1400 18700 1900 18700
rect 1400 18700 1900 18700
rect 1400 18700 1500 18700
rect 1800 18700 1900 18700
rect 1300 18700 1500 18800
rect 1800 18700 1900 18800
rect 1300 18800 1400 18800
rect 1800 18800 2000 18800
rect 1300 18800 1400 18800
rect 1900 18800 2000 18800
rect 1300 18800 1400 18800
rect 1900 18800 2000 18800
rect 1300 18800 1400 18800
rect 1900 18800 2000 18800
rect 1300 18800 1400 18900
rect 1900 18800 2000 18900
rect 1300 18900 1400 18900
rect 1900 18900 2000 18900
rect 1300 18900 1400 18900
rect 1900 18900 2000 18900
rect 1300 18900 1400 18900
rect 1900 18900 2000 18900
rect 1300 18900 1400 18900
rect 1900 18900 2000 18900
rect 1300 18900 1400 19000
rect 1900 18900 2000 19000
rect 1300 19000 1400 19000
rect 1900 19000 2000 19000
rect 1300 19000 1400 19000
rect 1900 19000 2000 19000
rect 1300 19000 1400 19000
rect 1900 19000 2000 19000
rect 1300 19000 1400 19000
rect 1900 19000 2000 19000
rect 1300 19000 1400 19100
rect 1900 19000 2000 19100
rect 1300 19100 1400 19100
rect 1800 19100 2000 19100
rect 1300 19100 1500 19100
rect 1800 19100 1900 19100
rect 1400 19100 1500 19100
rect 1700 19100 1900 19100
rect 1400 19100 1900 19100
rect 1400 19100 1900 19200
rect 1400 19200 1900 19200
rect 1500 19200 1800 19200
rect 1500 19200 1800 19200
rect 0 19700 500 19800
rect 0 19800 500 19800
rect 0 19800 500 19800
rect 0 19800 500 19800
rect 0 19800 500 19800
rect 0 19800 500 19900
rect 0 19900 500 19900
rect 0 19900 500 19900
rect 0 19900 500 19900
rect 0 19900 400 19900
rect 0 19900 400 20000
rect 0 20000 400 20000
rect 0 20000 400 20000
rect 0 20000 400 20000
rect 0 20000 400 20000
rect 0 20000 400 20100
rect 0 20100 400 20100
rect 0 20100 400 20100
rect 0 20100 300 20100
rect 0 20100 300 20100
rect 0 20100 300 20200
rect 0 20200 300 20200
rect 0 20200 200 20200
rect 0 20200 200 20200
rect 0 20200 200 20200
rect 0 20200 100 20300
rect 0 20300 100 20300
rect -600 0 -500 22000
rect 5500 0 5600 22000
<< labels >>
rlabel metal4 s 5500 0 5600 22000 6 vccd1
port 1 nsew power input
rlabel metal4 s -600 0 -500 22000 6 vssd1
port 2 nsew ground input
<< end >>
