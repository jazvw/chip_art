VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_art
  CLASS BLOCK ;
  FOREIGN chip_art ;
  ORIGIN 6.000 0.000 ;
  SIZE 62.000 BY 220.000 ;
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 55.000 0.000 56.000 220.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -6.000 0.000 -5.000 220.000 ;
    END
  END vssd1
  OBS
      LAYER met1 ;
        RECT 13.000 219.000 27.000 220.000 ;
        RECT 14.000 218.000 28.000 219.000 ;
        RECT 15.000 217.000 28.000 218.000 ;
        RECT 17.000 216.000 29.000 217.000 ;
        RECT 18.000 215.000 30.000 216.000 ;
        RECT 19.000 214.000 30.000 215.000 ;
        RECT 20.000 212.000 31.000 214.000 ;
        RECT 21.000 211.000 32.000 212.000 ;
        RECT 22.000 210.000 32.000 211.000 ;
        RECT 22.000 209.000 33.000 210.000 ;
        RECT 23.000 207.000 33.000 209.000 ;
        RECT 24.000 206.000 33.000 207.000 ;
        RECT 24.000 203.000 34.000 206.000 ;
        RECT 25.000 201.000 34.000 203.000 ;
        RECT 25.000 197.000 35.000 201.000 ;
        RECT 19.000 187.000 20.000 188.000 ;
        RECT 15.000 174.000 20.000 175.000 ;
        RECT 13.000 171.000 14.000 172.000 ;
        RECT 20.000 167.000 21.000 168.000 ;
        RECT 17.000 166.000 18.000 167.000 ;
        RECT 15.000 153.000 16.000 154.000 ;
        RECT 27.000 151.000 28.000 152.000 ;
        RECT 31.000 151.000 32.000 152.000 ;
        RECT 15.000 149.000 16.000 151.000 ;
        RECT 29.000 150.000 30.000 151.000 ;
        RECT 30.000 147.000 31.000 148.000 ;
        RECT 13.000 145.000 14.000 146.000 ;
        RECT 15.000 145.000 16.000 146.000 ;
        RECT 10.000 142.000 20.000 143.000 ;
        RECT 16.000 136.000 17.000 137.000 ;
        RECT 29.000 132.000 30.000 133.000 ;
        RECT 27.000 125.000 28.000 126.000 ;
        RECT 32.000 122.000 33.000 123.000 ;
        RECT 18.000 121.000 19.000 122.000 ;
        RECT 24.000 118.000 25.000 119.000 ;
        RECT 32.000 116.000 33.000 117.000 ;
        RECT 19.000 113.000 20.000 114.000 ;
        RECT 15.000 106.000 16.000 107.000 ;
        RECT 18.000 96.000 19.000 97.000 ;
        RECT 15.000 93.000 16.000 95.000 ;
        RECT 13.000 89.000 14.000 90.000 ;
        RECT 15.000 89.000 16.000 90.000 ;
        RECT 18.000 86.000 19.000 87.000 ;
        RECT 16.000 78.000 17.000 79.000 ;
        RECT 16.000 75.000 17.000 76.000 ;
        RECT 15.000 74.000 16.000 75.000 ;
        RECT 17.000 71.000 18.000 72.000 ;
        RECT 13.000 70.000 14.000 71.000 ;
      LAYER met2 ;
        RECT 0.000 219.000 13.000 220.000 ;
        RECT 0.000 218.000 14.000 219.000 ;
        RECT 0.000 217.000 15.000 218.000 ;
        RECT 0.000 216.000 17.000 217.000 ;
        RECT 0.000 215.000 18.000 216.000 ;
        RECT 0.000 214.000 19.000 215.000 ;
        RECT 0.000 213.000 20.000 214.000 ;
        RECT 3.000 212.000 20.000 213.000 ;
        RECT 6.000 211.000 21.000 212.000 ;
        RECT 8.000 210.000 22.000 211.000 ;
        RECT 9.000 209.000 22.000 210.000 ;
        RECT 10.000 208.000 23.000 209.000 ;
        RECT 11.000 207.000 23.000 208.000 ;
        RECT 12.000 206.000 24.000 207.000 ;
        RECT 13.000 204.000 24.000 206.000 ;
        RECT 14.000 203.000 24.000 204.000 ;
        RECT 14.000 201.000 25.000 203.000 ;
        RECT 15.000 197.000 25.000 201.000 ;
        RECT 18.000 190.000 19.000 191.000 ;
        RECT 14.000 186.000 15.000 187.000 ;
        RECT 13.000 152.000 14.000 153.000 ;
        RECT 27.000 152.000 28.000 153.000 ;
        RECT 16.000 150.000 17.000 151.000 ;
        RECT 13.000 149.000 14.000 150.000 ;
        RECT 10.000 141.000 14.000 142.000 ;
        RECT 16.000 141.000 17.000 142.000 ;
        RECT 19.000 141.000 20.000 142.000 ;
        RECT 26.000 141.000 27.000 142.000 ;
        RECT 25.000 135.000 26.000 136.000 ;
        RECT 31.000 135.000 32.000 136.000 ;
        RECT 30.000 130.000 31.000 131.000 ;
        RECT 13.000 129.000 14.000 130.000 ;
        RECT 27.000 121.000 28.000 122.000 ;
        RECT 30.000 121.000 31.000 122.000 ;
        RECT 18.000 116.000 19.000 117.000 ;
        RECT 14.000 112.000 15.000 113.000 ;
        RECT 16.000 108.000 17.000 110.000 ;
        RECT 15.000 105.000 16.000 106.000 ;
        RECT 16.000 94.000 17.000 95.000 ;
        RECT 13.000 93.000 14.000 94.000 ;
        RECT 13.000 71.000 14.000 72.000 ;
      LAYER met3 ;
        RECT 0.000 212.000 3.000 213.000 ;
        RECT 0.000 211.000 6.000 212.000 ;
        RECT 0.000 210.000 8.000 211.000 ;
        RECT 0.000 209.000 9.000 210.000 ;
        RECT 0.000 208.000 10.000 209.000 ;
        RECT 0.000 207.000 11.000 208.000 ;
        RECT 0.000 206.000 12.000 207.000 ;
        RECT 0.000 204.000 13.000 206.000 ;
        RECT 0.000 203.000 14.000 204.000 ;
        RECT 1.000 202.000 14.000 203.000 ;
        RECT 3.000 201.000 14.000 202.000 ;
        RECT 4.000 199.000 15.000 201.000 ;
        RECT 5.000 197.000 15.000 199.000 ;
      LAYER met4 ;
        RECT 0.000 202.000 1.000 203.000 ;
        RECT 0.000 201.000 3.000 202.000 ;
        RECT 0.000 199.000 4.000 201.000 ;
        RECT 0.000 197.000 5.000 199.000 ;
        RECT 14.000 191.000 19.000 192.000 ;
        RECT 13.000 188.000 14.000 191.000 ;
        RECT 19.000 188.000 20.000 191.000 ;
        RECT 13.000 187.000 15.000 188.000 ;
        RECT 18.000 187.000 19.000 188.000 ;
        RECT 15.000 186.000 18.000 187.000 ;
        RECT 13.000 183.000 14.000 185.000 ;
        RECT 19.000 183.000 20.000 185.000 ;
        RECT 11.000 182.000 19.000 183.000 ;
        RECT 13.000 181.000 14.000 182.000 ;
        RECT 15.000 175.000 20.000 176.000 ;
        RECT 13.000 174.000 15.000 175.000 ;
        RECT 13.000 172.000 14.000 174.000 ;
        RECT 13.000 170.000 20.000 171.000 ;
        RECT 13.000 167.000 20.000 168.000 ;
        RECT 14.000 166.000 15.000 167.000 ;
        RECT 18.000 166.000 19.000 167.000 ;
        RECT 20.000 166.000 22.000 167.000 ;
        RECT 13.000 163.000 14.000 166.000 ;
        RECT 19.000 164.000 20.000 166.000 ;
        RECT 18.000 163.000 20.000 164.000 ;
        RECT 21.000 163.000 22.000 166.000 ;
        RECT 14.000 162.000 19.000 163.000 ;
        RECT 10.000 159.000 12.000 160.000 ;
        RECT 13.000 159.000 20.000 160.000 ;
        RECT 13.000 153.000 14.000 157.000 ;
        RECT 17.000 156.000 19.000 157.000 ;
        RECT 23.000 156.000 29.000 157.000 ;
        RECT 30.000 156.000 32.000 157.000 ;
        RECT 16.000 153.000 17.000 156.000 ;
        RECT 14.000 152.000 16.000 153.000 ;
        RECT 19.000 152.000 20.000 156.000 ;
        RECT 25.000 152.000 27.000 153.000 ;
        RECT 28.000 151.000 31.000 152.000 ;
        RECT 30.000 150.000 32.000 151.000 ;
        RECT 14.000 149.000 15.000 150.000 ;
        RECT 13.000 146.000 14.000 149.000 ;
        RECT 16.000 146.000 17.000 150.000 ;
        RECT 19.000 146.000 20.000 150.000 ;
        RECT 26.000 149.000 29.000 150.000 ;
        RECT 25.000 148.000 27.000 149.000 ;
        RECT 27.000 147.000 30.000 148.000 ;
        RECT 30.000 146.000 32.000 147.000 ;
        RECT 14.000 145.000 15.000 146.000 ;
        RECT 16.000 145.000 19.000 146.000 ;
        RECT 26.000 145.000 30.000 146.000 ;
        RECT 15.000 144.000 18.000 145.000 ;
        RECT 25.000 144.000 26.000 145.000 ;
        RECT 25.000 142.000 27.000 143.000 ;
        RECT 14.000 141.000 16.000 142.000 ;
        RECT 17.000 141.000 19.000 142.000 ;
        RECT 27.000 141.000 29.000 142.000 ;
        RECT 13.000 138.000 14.000 141.000 ;
        RECT 19.000 138.000 20.000 141.000 ;
        RECT 29.000 140.000 32.000 141.000 ;
        RECT 30.000 139.000 32.000 140.000 ;
        RECT 27.000 138.000 30.000 139.000 ;
        RECT 14.000 137.000 19.000 138.000 ;
        RECT 25.000 137.000 27.000 138.000 ;
        RECT 25.000 134.000 27.000 135.000 ;
        RECT 13.000 130.000 14.000 132.000 ;
        RECT 25.000 130.000 26.000 134.000 ;
        RECT 27.000 133.000 28.000 134.000 ;
        RECT 28.000 132.000 29.000 133.000 ;
        RECT 31.000 132.000 32.000 135.000 ;
        RECT 29.000 131.000 32.000 132.000 ;
        RECT 31.000 130.000 32.000 131.000 ;
        RECT 13.000 128.000 20.000 129.000 ;
        RECT 22.000 127.000 24.000 128.000 ;
        RECT 25.000 127.000 34.000 128.000 ;
        RECT 33.000 126.000 34.000 127.000 ;
        RECT 13.000 125.000 20.000 126.000 ;
        RECT 18.000 124.000 19.000 125.000 ;
        RECT 25.000 124.000 27.000 125.000 ;
        RECT 29.000 124.000 30.000 125.000 ;
        RECT 19.000 121.000 20.000 124.000 ;
        RECT 24.000 122.000 25.000 124.000 ;
        RECT 30.000 123.000 31.000 124.000 ;
        RECT 32.000 123.000 33.000 124.000 ;
        RECT 26.000 122.000 31.000 123.000 ;
        RECT 13.000 120.000 19.000 121.000 ;
        RECT 23.000 119.000 24.000 122.000 ;
        RECT 26.000 119.000 27.000 121.000 ;
        RECT 30.000 119.000 31.000 121.000 ;
        RECT 27.000 118.000 31.000 119.000 ;
        RECT 33.000 118.000 34.000 122.000 ;
        RECT 14.000 117.000 19.000 118.000 ;
        RECT 24.000 117.000 25.000 118.000 ;
        RECT 32.000 117.000 33.000 118.000 ;
        RECT 13.000 114.000 14.000 117.000 ;
        RECT 19.000 114.000 20.000 117.000 ;
        RECT 25.000 116.000 26.000 117.000 ;
        RECT 31.000 116.000 32.000 117.000 ;
        RECT 26.000 115.000 31.000 116.000 ;
        RECT 13.000 113.000 15.000 114.000 ;
        RECT 18.000 113.000 19.000 114.000 ;
        RECT 15.000 112.000 18.000 113.000 ;
        RECT 13.000 110.000 14.000 111.000 ;
        RECT 14.000 109.000 16.000 110.000 ;
        RECT 17.000 108.000 19.000 109.000 ;
        RECT 18.000 107.000 21.000 108.000 ;
        RECT 16.000 106.000 18.000 107.000 ;
        RECT 13.000 105.000 15.000 106.000 ;
        RECT 21.000 105.000 22.000 107.000 ;
        RECT 13.000 97.000 14.000 100.000 ;
        RECT 19.000 98.000 20.000 100.000 ;
        RECT 18.000 97.000 20.000 98.000 ;
        RECT 11.000 96.000 18.000 97.000 ;
        RECT 14.000 93.000 15.000 94.000 ;
        RECT 13.000 90.000 14.000 93.000 ;
        RECT 16.000 90.000 17.000 94.000 ;
        RECT 19.000 90.000 20.000 94.000 ;
        RECT 14.000 89.000 15.000 90.000 ;
        RECT 16.000 89.000 19.000 90.000 ;
        RECT 15.000 88.000 18.000 89.000 ;
        RECT 14.000 86.000 17.000 87.000 ;
        RECT 13.000 82.000 14.000 86.000 ;
        RECT 16.000 82.000 17.000 86.000 ;
        RECT 19.000 83.000 20.000 86.000 ;
        RECT 18.000 82.000 20.000 83.000 ;
        RECT 14.000 81.000 19.000 82.000 ;
        RECT 13.000 78.000 16.000 79.000 ;
        RECT 16.000 77.000 20.000 78.000 ;
        RECT 17.000 76.000 20.000 77.000 ;
        RECT 13.000 75.000 16.000 76.000 ;
        RECT 13.000 74.000 15.000 75.000 ;
        RECT 16.000 73.000 19.000 74.000 ;
        RECT 17.000 72.000 20.000 73.000 ;
        RECT 11.000 69.000 12.000 72.000 ;
        RECT 14.000 71.000 17.000 72.000 ;
        RECT 11.000 67.000 20.000 69.000 ;
        RECT 11.000 64.000 12.000 67.000 ;
        RECT 21.000 55.000 28.000 56.000 ;
        RECT 17.000 54.000 32.000 55.000 ;
        RECT 14.000 53.000 35.000 54.000 ;
        RECT 12.000 52.000 37.000 53.000 ;
        RECT 11.000 51.000 38.000 52.000 ;
        RECT 10.000 50.000 40.000 51.000 ;
        RECT 8.000 49.000 41.000 50.000 ;
        RECT 7.000 48.000 42.000 49.000 ;
        RECT 6.000 47.000 43.000 48.000 ;
        RECT 6.000 46.000 44.000 47.000 ;
        RECT 5.000 45.000 44.000 46.000 ;
        RECT 4.000 44.000 45.000 45.000 ;
        RECT 4.000 43.000 15.000 44.000 ;
        RECT 17.000 43.000 33.000 44.000 ;
        RECT 34.000 43.000 46.000 44.000 ;
        RECT 3.000 42.000 13.000 43.000 ;
        RECT 19.000 42.000 30.000 43.000 ;
        RECT 36.000 42.000 46.000 43.000 ;
        RECT 3.000 41.000 12.000 42.000 ;
        RECT 2.000 39.000 12.000 41.000 ;
        RECT 1.000 37.000 12.000 39.000 ;
        RECT 20.000 37.000 29.000 42.000 ;
        RECT 37.000 40.000 47.000 42.000 ;
        RECT 38.000 39.000 47.000 40.000 ;
        RECT 1.000 36.000 13.000 37.000 ;
        RECT 19.000 36.000 30.000 37.000 ;
        RECT 37.000 36.000 48.000 39.000 ;
        RECT 1.000 35.000 14.000 36.000 ;
        RECT 18.000 35.000 31.000 36.000 ;
        RECT 35.000 35.000 48.000 36.000 ;
        RECT 1.000 33.000 48.000 35.000 ;
        RECT 1.000 30.000 49.000 33.000 ;
        RECT 1.000 29.000 12.000 30.000 ;
        RECT 13.000 29.000 35.000 30.000 ;
        RECT 1.000 25.000 10.000 29.000 ;
        RECT 14.000 27.000 35.000 29.000 ;
        RECT 14.000 26.000 34.000 27.000 ;
        RECT 15.000 25.000 34.000 26.000 ;
        RECT 39.000 25.000 48.000 30.000 ;
        RECT 2.000 23.000 11.000 25.000 ;
        RECT 16.000 24.000 33.000 25.000 ;
        RECT 16.000 23.000 32.000 24.000 ;
        RECT 38.000 23.000 47.000 25.000 ;
        RECT 2.000 22.000 12.000 23.000 ;
        RECT 18.000 22.000 31.000 23.000 ;
        RECT 37.000 22.000 47.000 23.000 ;
        RECT 3.000 21.000 13.000 22.000 ;
        RECT 19.000 21.000 30.000 22.000 ;
        RECT 36.000 21.000 46.000 22.000 ;
        RECT 3.000 20.000 14.000 21.000 ;
        RECT 22.000 20.000 27.000 21.000 ;
        RECT 35.000 20.000 46.000 21.000 ;
        RECT 4.000 19.000 15.000 20.000 ;
        RECT 34.000 19.000 45.000 20.000 ;
        RECT 4.000 18.000 16.000 19.000 ;
        RECT 33.000 18.000 45.000 19.000 ;
        RECT 5.000 17.000 18.000 18.000 ;
        RECT 31.000 17.000 44.000 18.000 ;
        RECT 6.000 16.000 20.000 17.000 ;
        RECT 29.000 16.000 43.000 17.000 ;
        RECT 7.000 15.000 42.000 16.000 ;
        RECT 8.000 14.000 41.000 15.000 ;
        RECT 9.000 13.000 40.000 14.000 ;
        RECT 10.000 12.000 39.000 13.000 ;
        RECT 12.000 11.000 38.000 12.000 ;
        RECT 13.000 10.000 36.000 11.000 ;
        RECT 15.000 9.000 34.000 10.000 ;
        RECT 18.000 8.000 31.000 9.000 ;
  END
END chip_art
END LIBRARY

