/* SPDX-FileCopyrightText: 2022 Jasper van Woudenberg
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0
*/


// This is here to keep various parts of the hardening flow happy
module chip_art(
`ifdef USE_POWER_PINS
        input vccd1,
        input vssd1,
`endif
        input wb_clk_i,
        input active

);
endmodule
