../../gds/chip_art.lef